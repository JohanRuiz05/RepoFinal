* NGSPICE file created from tt_um_mult_4.ext - technology: sky130A

X0 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=2.48945k ps=24.76584k w=0.87 l=1.97
X1 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=1.5774k ps=17.7898k w=0.55 l=1.97
X2 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X13 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X14 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X15 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X16 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X17 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X18 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X19 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X20 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X21 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X22 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X23 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X24 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X25 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X26 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X27 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X28 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X29 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X30 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X31 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X32 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X33 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X34 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X35 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X36 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X37 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X38 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X39 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X40 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X41 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X42 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X43 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X44 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X45 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X46 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X47 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X48 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X49 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X50 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X51 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X52 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X53 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X54 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X55 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X56 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X57 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X58 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X59 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X60 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X61 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X62 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X63 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X64 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X65 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X66 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X67 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X68 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X69 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X70 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X71 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X72 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X73 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X74 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X75 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X76 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X77 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X78 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X79 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X80 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X81 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X82 uo_out[6] _277_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X83 _277_/a_1020_47# _277_/a_27_47# _277_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X84 _277_/a_572_47# _277_/a_193_47# _277_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X85 VPWR _277_/a_1062_300# _277_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X86 _277_/a_634_183# _277_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X87 VPWR _277_/CLK _277_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X88 _277_/a_381_47# _277_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X89 _277_/a_475_413# _277_/a_27_47# _277_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X90 VGND _277_/a_1062_300# _277_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X91 VPWR _277_/a_634_183# _277_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X92 uo_out[6] _277_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09262 ps=0.935 w=0.65 l=0.15
X93 _277_/a_568_413# _277_/a_27_47# _277_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X94 _277_/a_634_183# _277_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X95 _277_/a_975_413# _277_/a_193_47# _277_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X96 _277_/a_193_47# _277_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X97 _277_/a_891_413# _277_/a_27_47# _277_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X98 uo_out[6] _277_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10563 ps=0.975 w=0.65 l=0.15
X99 VGND _277_/a_891_413# _277_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X100 VPWR _277_/a_1062_300# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X101 VGND _277_/a_1062_300# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X102 uo_out[6] _277_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X103 _277_/a_193_47# _277_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X104 VGND _277_/a_1062_300# uo_out[6] VGND sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 _277_/a_381_47# _277_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X106 VPWR _277_/a_891_413# _277_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X107 _277_/a_475_413# _277_/a_193_47# _277_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X108 _277_/a_891_413# _277_/a_193_47# _277_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X109 VGND _277_/a_634_183# _277_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X110 VGND _277_/CLK _277_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X111 VPWR _277_/a_1062_300# uo_out[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X148 VGND _256_/Q _200_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X149 _200_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X150 _200_/X _200_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X151 VPWR _256_/Q _200_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X152 _200_/X _200_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X153 _200_/a_150_297# _202_/B _200_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X158 _131_/Y _133_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X159 VGND _133_/A _131_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X160 _131_/Y _133_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 VPWR _133_/A _131_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X400 _264_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X401 VGND _285_/CLK _264_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X402 _264_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X403 VPWR _285_/CLK _264_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X418 uo_out[5] _276_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X419 _276_/a_1020_47# _276_/a_27_47# _276_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X420 _276_/a_572_47# _276_/a_193_47# _276_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X421 VPWR _276_/a_1062_300# _276_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X422 _276_/a_634_183# _276_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X423 VPWR _276_/CLK _276_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X424 _276_/a_381_47# _276_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X425 _276_/a_475_413# _276_/a_27_47# _276_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X426 VGND _276_/a_1062_300# _276_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X427 VPWR _276_/a_634_183# _276_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X428 uo_out[5] _276_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X429 _276_/a_568_413# _276_/a_27_47# _276_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X430 _276_/a_634_183# _276_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X431 _276_/a_975_413# _276_/a_193_47# _276_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X432 _276_/a_193_47# _276_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X433 _276_/a_891_413# _276_/a_27_47# _276_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X434 uo_out[5] _276_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X435 VGND _276_/a_891_413# _276_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X436 VPWR _276_/a_1062_300# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X437 VGND _276_/a_1062_300# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X438 uo_out[5] _276_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 _276_/a_193_47# _276_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X440 VGND _276_/a_1062_300# uo_out[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X441 _276_/a_381_47# _276_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X442 VPWR _276_/a_891_413# _276_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X443 _276_/a_475_413# _276_/a_193_47# _276_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X444 _276_/a_891_413# _276_/a_193_47# _276_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X445 VGND _276_/a_634_183# _276_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X446 VGND _276_/CLK _276_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X447 VPWR _276_/a_1062_300# uo_out[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X482 VPWR uo_out[6] _133_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X483 _133_/A uo_out[6] _130_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X484 _130_/a_113_47# _260_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X485 _133_/A _260_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X504 hold8/A _259_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X505 _259_/a_891_413# _259_/a_193_47# _259_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X506 _259_/a_561_413# _259_/a_27_47# _259_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X507 VPWR _259_/CLK _259_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X508 hold8/A _259_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X509 _259_/a_381_47# _259_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X510 VGND _259_/a_634_159# _259_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X511 VPWR _259_/a_891_413# _259_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X512 _259_/a_466_413# _259_/a_193_47# _259_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X513 VPWR _259_/a_634_159# _259_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X514 _259_/a_634_159# _259_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X515 _259_/a_634_159# _259_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X516 _259_/a_975_413# _259_/a_193_47# _259_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X517 VGND _259_/a_1059_315# _259_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X518 _259_/a_193_47# _259_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X519 _259_/a_891_413# _259_/a_27_47# _259_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X520 _259_/a_592_47# _259_/a_193_47# _259_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X521 VPWR _259_/a_1059_315# _259_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X522 _259_/a_1017_47# _259_/a_27_47# _259_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X523 _259_/a_193_47# _259_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X524 _259_/a_466_413# _259_/a_27_47# _259_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X525 VGND _259_/a_891_413# _259_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X526 _259_/a_381_47# _259_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X527 VGND _259_/CLK _259_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X596 VPWR _263_/Q hold20/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X597 VGND hold20/a_285_47# hold20/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X598 hold20/X hold20/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X599 VGND _263_/Q hold20/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X600 VPWR hold20/a_285_47# hold20/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X601 hold20/a_285_47# hold20/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X602 hold20/a_285_47# hold20/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X603 hold20/X hold20/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X770 uo_out[4] _275_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X771 _275_/a_1020_47# _275_/a_27_47# _275_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X772 _275_/a_572_47# _275_/a_193_47# _275_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X773 VPWR _275_/a_1062_300# _275_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X774 _275_/a_634_183# _275_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X775 VPWR _275_/CLK _275_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X776 _275_/a_381_47# _275_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X777 _275_/a_475_413# _275_/a_27_47# _275_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X778 VGND _275_/a_1062_300# _275_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X779 VPWR _275_/a_634_183# _275_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X780 uo_out[4] _275_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X781 _275_/a_568_413# _275_/a_27_47# _275_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X782 _275_/a_634_183# _275_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X783 _275_/a_975_413# _275_/a_193_47# _275_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X784 _275_/a_193_47# _275_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X785 _275_/a_891_413# _275_/a_27_47# _275_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X786 uo_out[4] _275_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X787 VGND _275_/a_891_413# _275_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X788 VPWR _275_/a_1062_300# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X789 VGND _275_/a_1062_300# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X790 uo_out[4] _275_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X791 _275_/a_193_47# _275_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X792 VGND _275_/a_1062_300# uo_out[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X793 _275_/a_381_47# _275_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X794 VPWR _275_/a_891_413# _275_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X795 _275_/a_475_413# _275_/a_193_47# _275_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X796 _275_/a_891_413# _275_/a_193_47# _275_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X797 VGND _275_/a_634_183# _275_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X798 VGND _275_/CLK _275_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X799 VPWR _275_/a_1062_300# uo_out[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X858 _258_/Q _258_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X859 _258_/a_891_413# _258_/a_193_47# _258_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X860 _258_/a_561_413# _258_/a_27_47# _258_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X861 VPWR _258_/CLK _258_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X862 _258_/Q _258_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X863 _258_/a_381_47# _258_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X864 VGND _258_/a_634_159# _258_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X865 VPWR _258_/a_891_413# _258_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X866 _258_/a_466_413# _258_/a_193_47# _258_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X867 VPWR _258_/a_634_159# _258_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X868 _258_/a_634_159# _258_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X869 _258_/a_634_159# _258_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X870 _258_/a_975_413# _258_/a_193_47# _258_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X871 VGND _258_/a_1059_315# _258_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X872 _258_/a_193_47# _258_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X873 _258_/a_891_413# _258_/a_27_47# _258_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X874 _258_/a_592_47# _258_/a_193_47# _258_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X875 VPWR _258_/a_1059_315# _258_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X876 _258_/a_1017_47# _258_/a_27_47# _258_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X877 _258_/a_193_47# _258_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X878 _258_/a_466_413# _258_/a_27_47# _258_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X879 VGND _258_/a_891_413# _258_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X880 _258_/a_381_47# _258_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X881 VGND _258_/CLK _258_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X882 _189_/a_240_47# input7/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X883 _265_/D _189_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X884 VGND _203_/A1 _189_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X885 _189_/a_51_297# hold6/X _189_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X886 _189_/a_149_47# _188_/X _189_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X887 _189_/a_240_47# _186_/Y _189_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X888 VPWR _203_/A1 _189_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X889 _265_/D _189_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X890 _189_/a_149_47# hold6/X _189_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X891 _189_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X892 VPWR _188_/X _189_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X893 _189_/a_512_297# input7/X _189_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X970 VPWR _268_/Q hold10/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X971 VGND hold10/a_285_47# hold10/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X972 hold10/X hold10/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X973 VGND _268_/Q hold10/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X974 VPWR hold10/a_285_47# hold10/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X975 hold10/a_285_47# hold10/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X976 hold10/a_285_47# hold10/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X977 hold10/X hold10/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1148 uo_out[3] _274_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X1149 _274_/a_1020_47# _274_/a_27_47# _274_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X1150 _274_/a_572_47# _274_/a_193_47# _274_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X1151 VPWR _274_/a_1062_300# _274_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X1152 _274_/a_634_183# _274_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X1153 VPWR _274_/CLK _274_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1154 _274_/a_381_47# _274_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X1155 _274_/a_475_413# _274_/a_27_47# _274_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X1156 VGND _274_/a_1062_300# _274_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1157 VPWR _274_/a_634_183# _274_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1158 uo_out[3] _274_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1159 _274_/a_568_413# _274_/a_27_47# _274_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X1160 _274_/a_634_183# _274_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1161 _274_/a_975_413# _274_/a_193_47# _274_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1162 _274_/a_193_47# _274_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1163 _274_/a_891_413# _274_/a_27_47# _274_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1164 uo_out[3] _274_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1165 VGND _274_/a_891_413# _274_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1166 VPWR _274_/a_1062_300# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1167 VGND _274_/a_1062_300# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1168 uo_out[3] _274_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1169 _274_/a_193_47# _274_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1170 VGND _274_/a_1062_300# uo_out[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1171 _274_/a_381_47# _274_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1172 VPWR _274_/a_891_413# _274_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X1173 _274_/a_475_413# _274_/a_193_47# _274_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1174 _274_/a_891_413# _274_/a_193_47# _274_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1175 VGND _274_/a_634_183# _274_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1176 VGND _274_/CLK _274_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1177 VPWR _274_/a_1062_300# uo_out[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1180 _260_/CLK _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1181 VGND _267_/CLK _260_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1182 _260_/CLK _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1183 VPWR _267_/CLK _260_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1244 _257_/Q _257_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1245 _257_/a_891_413# _257_/a_193_47# _257_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1246 _257_/a_561_413# _257_/a_27_47# _257_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1247 VPWR _257_/CLK _257_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1248 _257_/Q _257_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1249 _257_/a_381_47# _257_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1250 VGND _257_/a_634_159# _257_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1251 VPWR _257_/a_891_413# _257_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1252 _257_/a_466_413# _257_/a_193_47# _257_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1253 VPWR _257_/a_634_159# _257_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1254 _257_/a_634_159# _257_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1255 _257_/a_634_159# _257_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1256 _257_/a_975_413# _257_/a_193_47# _257_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1257 VGND _257_/a_1059_315# _257_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1258 _257_/a_193_47# _257_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1259 _257_/a_891_413# _257_/a_27_47# _257_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1260 _257_/a_592_47# _257_/a_193_47# _257_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1261 VPWR _257_/a_1059_315# _257_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1262 _257_/a_1017_47# _257_/a_27_47# _257_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1263 _257_/a_193_47# _257_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1264 _257_/a_466_413# _257_/a_27_47# _257_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1265 VGND _257_/a_891_413# _257_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1266 _257_/a_381_47# _257_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1267 VGND _257_/CLK _257_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1268 VGND _265_/Q _188_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1269 _188_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1270 _188_/X _188_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1271 VPWR _265_/Q _188_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1272 _188_/X _188_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1273 _188_/a_150_297# _202_/B _188_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1358 VPWR _265_/Q hold11/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1359 VGND hold11/a_285_47# hold11/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1360 hold11/X hold11/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1361 VGND _265_/Q hold11/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1362 VPWR hold11/a_285_47# hold11/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1363 hold11/a_285_47# hold11/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1364 hold11/a_285_47# hold11/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1365 hold11/X hold11/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1506 uo_out[2] _273_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X1507 _273_/a_1020_47# _273_/a_27_47# _273_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X1508 _273_/a_572_47# _273_/a_193_47# _273_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X1509 VPWR _273_/a_1062_300# _273_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X1510 _273_/a_634_183# _273_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X1511 VPWR _273_/CLK _273_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1512 _273_/a_381_47# _273_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X1513 _273_/a_475_413# _273_/a_27_47# _273_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X1514 VGND _273_/a_1062_300# _273_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1515 VPWR _273_/a_634_183# _273_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1516 uo_out[2] _273_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1517 _273_/a_568_413# _273_/a_27_47# _273_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X1518 _273_/a_634_183# _273_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1519 _273_/a_975_413# _273_/a_193_47# _273_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1520 _273_/a_193_47# _273_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1521 _273_/a_891_413# _273_/a_27_47# _273_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1522 uo_out[2] _273_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1523 VGND _273_/a_891_413# _273_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1524 VPWR _273_/a_1062_300# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1525 VGND _273_/a_1062_300# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1526 uo_out[2] _273_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1527 _273_/a_193_47# _273_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1528 VGND _273_/a_1062_300# uo_out[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1529 _273_/a_381_47# _273_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1530 VPWR _273_/a_891_413# _273_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X1531 _273_/a_475_413# _273_/a_193_47# _273_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1532 _273_/a_891_413# _273_/a_193_47# _273_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1533 VGND _273_/a_634_183# _273_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1534 VGND _273_/CLK _273_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1535 VPWR _273_/a_1062_300# uo_out[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1596 _256_/Q _256_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1597 _256_/a_891_413# _256_/a_193_47# _256_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1598 _256_/a_561_413# _256_/a_27_47# _256_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1599 VPWR _256_/CLK _256_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1600 _256_/Q _256_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1601 _256_/a_381_47# _256_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1602 VGND _256_/a_634_159# _256_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1603 VPWR _256_/a_891_413# _256_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1604 _256_/a_466_413# _256_/a_193_47# _256_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1605 VPWR _256_/a_634_159# _256_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1606 _256_/a_634_159# _256_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1607 _256_/a_634_159# _256_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1608 _256_/a_975_413# _256_/a_193_47# _256_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1609 VGND _256_/a_1059_315# _256_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1610 _256_/a_193_47# _256_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1611 _256_/a_891_413# _256_/a_27_47# _256_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1612 _256_/a_592_47# _256_/a_193_47# _256_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1613 VPWR _256_/a_1059_315# _256_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1614 _256_/a_1017_47# _256_/a_27_47# _256_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1615 _256_/a_193_47# _256_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1616 _256_/a_466_413# _256_/a_27_47# _256_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1617 VGND _256_/a_891_413# _256_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 _256_/a_381_47# _256_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1619 VGND _256_/CLK _256_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1620 _187_/a_240_47# input8/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1621 _266_/D _187_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1622 VGND _186_/A _187_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1623 _187_/a_51_297# hold1/X _187_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1624 _187_/a_149_47# _184_/X _187_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1625 _187_/a_240_47# _186_/Y _187_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1626 VPWR _186_/A _187_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1627 _266_/D _187_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1628 _187_/a_149_47# hold1/X _187_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1629 _187_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1630 VPWR _184_/X _187_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1631 _187_/a_512_297# input8/X _187_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1632 _262_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1633 VGND _285_/CLK _262_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1634 _262_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1635 VPWR _285_/CLK _262_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1662 clkload0/Y _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1663 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1664 clkload0/Y _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1665 clkload0/Y _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1667 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X1668 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1669 clkload0/Y _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1670 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1671 VGND _267_/CLK clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1672 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X1673 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1674 VGND _267_/CLK clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1675 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1676 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1677 VGND _267_/CLK clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1678 VPWR _267_/CLK clkload0/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1679 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1680 clkload0/Y _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1681 VGND _267_/CLK clkload0/Y VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1722 VPWR _258_/Q hold12/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1723 VGND hold12/a_285_47# hold12/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1724 hold12/X hold12/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1725 VGND _258_/Q hold12/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1726 VPWR hold12/a_285_47# hold12/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1727 hold12/a_285_47# hold12/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1728 hold12/a_285_47# hold12/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1729 hold12/X hold12/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1896 uo_out[1] _272_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X1897 _272_/a_1020_47# _272_/a_27_47# _272_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X1898 _272_/a_572_47# _272_/a_193_47# _272_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X1899 VPWR _272_/a_1062_300# _272_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X1900 _272_/a_634_183# _272_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X1901 VPWR _272_/CLK _272_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1902 _272_/a_381_47# _272_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X1903 _272_/a_475_413# _272_/a_27_47# _272_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X1904 VGND _272_/a_1062_300# _272_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1905 VPWR _272_/a_634_183# _272_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1906 uo_out[1] _272_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1907 _272_/a_568_413# _272_/a_27_47# _272_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X1908 _272_/a_634_183# _272_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1909 _272_/a_975_413# _272_/a_193_47# _272_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1910 _272_/a_193_47# _272_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1911 _272_/a_891_413# _272_/a_27_47# _272_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1912 uo_out[1] _272_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1913 VGND _272_/a_891_413# _272_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1914 VPWR _272_/a_1062_300# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1915 VGND _272_/a_1062_300# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1916 uo_out[1] _272_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1917 _272_/a_193_47# _272_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1918 VGND _272_/a_1062_300# uo_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1919 _272_/a_381_47# _272_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1920 VPWR _272_/a_891_413# _272_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X1921 _272_/a_475_413# _272_/a_193_47# _272_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1922 _272_/a_891_413# _272_/a_193_47# _272_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1923 VGND _272_/a_634_183# _272_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1924 VGND _272_/CLK _272_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1925 VPWR _272_/a_1062_300# uo_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1992 _255_/Q _255_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1993 _255_/a_891_413# _255_/a_193_47# _255_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1994 _255_/a_561_413# _255_/a_27_47# _255_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1995 VPWR _255_/CLK _255_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1996 _255_/Q _255_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1997 _255_/a_381_47# _255_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1998 VGND _255_/a_634_159# _255_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1999 VPWR _255_/a_891_413# _255_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2000 _255_/a_466_413# _255_/a_193_47# _255_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2001 VPWR _255_/a_634_159# _255_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2002 _255_/a_634_159# _255_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2003 _255_/a_634_159# _255_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2004 _255_/a_975_413# _255_/a_193_47# _255_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2005 VGND _255_/a_1059_315# _255_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2006 _255_/a_193_47# _255_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2007 _255_/a_891_413# _255_/a_27_47# _255_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2008 _255_/a_592_47# _255_/a_193_47# _255_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2009 VPWR _255_/a_1059_315# _255_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2010 _255_/a_1017_47# _255_/a_27_47# _255_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2011 _255_/a_193_47# _255_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2012 _255_/a_466_413# _255_/a_27_47# _255_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2013 VGND _255_/a_891_413# _255_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2014 _255_/a_381_47# _255_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2015 VGND _255_/CLK _255_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2020 VPWR _186_/A _186_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2021 _186_/Y _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2022 VPWR _269_/Q _186_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2023 _186_/a_27_47# _269_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2024 _186_/a_27_47# _186_/A _186_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2025 _186_/Y _186_/A _186_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2026 _186_/Y _269_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2027 VGND _269_/Q _186_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2058 VPWR clkload1/A clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2059 clkload1/Y clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2060 clkload1/Y clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2061 VPWR clkload1/A clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2062 clkload1/Y clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2063 VPWR clkload1/A clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2064 clkload1/Y clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X2065 clkload1/Y clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2066 clkload1/Y clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X2067 VGND clkload1/A clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2068 VGND clkload1/A clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2069 VGND clkload1/A clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X2070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2096 VGND _178_/A _169_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2097 _169_/a_510_47# _168_/X _169_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2098 _169_/a_79_21# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X2099 VPWR _168_/X _169_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X2100 _169_/a_79_21# uo_out[4] _169_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X2101 _169_/a_297_297# _178_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2102 _169_/a_79_21# _186_/A _169_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X2103 VPWR _169_/a_79_21# _275_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2104 VGND _169_/a_79_21# _275_/D VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2105 _169_/a_215_47# uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
X2106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2130 VPWR _301_/A hold13/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2131 VGND hold13/a_285_47# hold13/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2132 hold13/X hold13/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2133 VGND _301_/A hold13/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2134 VPWR hold13/a_285_47# hold13/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2135 hold13/a_285_47# hold13/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2136 hold13/a_285_47# hold13/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2137 hold13/X hold13/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2172 VPWR tt_um_mult_4_20/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2173 uio_oe[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2282 uo_out[0] _271_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2283 VPWR _271_/a_1059_315# uo_out[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2284 _271_/a_891_413# _271_/a_193_47# _271_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2285 _271_/a_561_413# _271_/a_27_47# _271_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2286 VPWR _271_/CLK _271_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2287 uo_out[0] _271_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2288 _271_/a_381_47# _271_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2289 VGND _271_/a_634_159# _271_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2290 VGND _271_/a_1059_315# uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2291 VPWR _271_/a_891_413# _271_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2292 _271_/a_466_413# _271_/a_193_47# _271_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2293 VPWR _271_/a_634_159# _271_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2294 _271_/a_634_159# _271_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2295 _271_/a_634_159# _271_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X2296 _271_/a_975_413# _271_/a_193_47# _271_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2297 VGND _271_/a_1059_315# _271_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2298 _271_/a_193_47# _271_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2299 _271_/a_891_413# _271_/a_27_47# _271_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2300 _271_/a_592_47# _271_/a_193_47# _271_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2301 VPWR _271_/a_1059_315# _271_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2302 _271_/a_1017_47# _271_/a_27_47# _271_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2303 _271_/a_193_47# _271_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2304 _271_/a_466_413# _271_/a_27_47# _271_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2305 VGND _271_/a_891_413# _271_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2306 _271_/a_381_47# _271_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2307 VGND _271_/CLK _271_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2370 _254_/Q _254_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2371 _254_/a_891_413# _254_/a_193_47# _254_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2372 _254_/a_561_413# _254_/a_27_47# _254_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2373 VPWR _254_/CLK _254_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2374 _254_/Q _254_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2375 _254_/a_381_47# _254_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2376 VGND _254_/a_634_159# _254_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2377 VPWR _254_/a_891_413# _254_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2378 _254_/a_466_413# _254_/a_193_47# _254_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2379 VPWR _254_/a_634_159# _254_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2380 _254_/a_634_159# _254_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2381 _254_/a_634_159# _254_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2382 _254_/a_975_413# _254_/a_193_47# _254_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2383 VGND _254_/a_1059_315# _254_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2384 _254_/a_193_47# _254_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2385 _254_/a_891_413# _254_/a_27_47# _254_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2386 _254_/a_592_47# _254_/a_193_47# _254_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2387 VPWR _254_/a_1059_315# _254_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2388 _254_/a_1017_47# _254_/a_27_47# _254_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2389 _254_/a_193_47# _254_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2390 _254_/a_466_413# _254_/a_27_47# _254_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2391 VGND _254_/a_891_413# _254_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2392 _254_/a_381_47# _254_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2393 VGND _254_/CLK _254_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2396 VPWR _269_/Q _185_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2397 _185_/X _185_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2398 VGND _269_/Q _185_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2399 _185_/a_59_75# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2400 _185_/X _185_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X2401 _185_/a_145_75# _186_/A _185_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2440 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2442 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2443 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X2444 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2445 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2446 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2447 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2448 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2449 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2450 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2451 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X2452 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2453 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2454 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2455 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2456 clkload2/Y _284_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2457 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2458 VPWR _284_/CLK clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2459 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2460 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2461 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2462 clkload2/Y _284_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2463 VGND _284_/CLK clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2480 _168_/a_81_21# _128_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X2481 _168_/a_299_297# _128_/Y _168_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2482 VPWR _168_/a_81_21# _168_/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2483 VPWR _151_/Y _168_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2484 VGND _168_/a_81_21# _168_/X VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2485 VGND _167_/X _168_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2486 _168_/a_299_297# _167_/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2487 _168_/a_384_47# _151_/Y _168_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X2488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2504 VPWR _279_/Q hold14/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2505 VGND hold14/a_285_47# hold14/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2506 _216_/A hold14/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2507 VGND _279_/Q hold14/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2508 VPWR hold14/a_285_47# hold14/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2509 hold14/a_285_47# hold14/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2510 hold14/a_285_47# hold14/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2511 _216_/A hold14/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2546 VPWR tt_um_mult_4_21/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2547 uio_oe[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2612 _271_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2613 VGND clkload1/A _271_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2614 _271_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2615 VPWR clkload1/A _271_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2656 _270_/Q _270_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2657 _270_/a_891_413# _270_/a_193_47# _270_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2658 _270_/a_561_413# _270_/a_27_47# _270_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2659 VPWR _284_/CLK _270_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2660 _270_/Q _270_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2661 _270_/a_381_47# _270_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2662 VGND _270_/a_634_159# _270_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2663 VPWR _270_/a_891_413# _270_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2664 _270_/a_466_413# _270_/a_193_47# _270_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2665 VPWR _270_/a_634_159# _270_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2666 _270_/a_634_159# _270_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2667 _270_/a_634_159# _270_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2668 _270_/a_975_413# _270_/a_193_47# _270_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2669 VGND _270_/a_1059_315# _270_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2670 _270_/a_193_47# _270_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2671 _270_/a_891_413# _270_/a_27_47# _270_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2672 _270_/a_592_47# _270_/a_193_47# _270_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2673 VPWR _270_/a_1059_315# _270_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2674 _270_/a_1017_47# _270_/a_27_47# _270_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2675 _270_/a_193_47# _270_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2676 _270_/a_466_413# _270_/a_27_47# _270_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2677 VGND _270_/a_891_413# _270_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2678 _270_/a_381_47# _270_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2679 VGND _284_/CLK _270_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2728 VGND hold7/X _184_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2729 _184_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2730 _184_/X _184_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2731 VPWR hold7/X _184_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2732 _184_/X _184_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2733 _184_/a_150_297# _202_/B _184_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2796 _167_/a_81_21# _151_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2797 _167_/a_299_297# _151_/A _167_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2798 VPWR _167_/a_81_21# _167_/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2799 VPWR _171_/B _167_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2800 VGND _167_/a_81_21# _167_/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2801 VGND _151_/C _167_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2802 _167_/a_299_297# _151_/C VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2803 _167_/a_384_47# _171_/B _167_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2820 VPWR _257_/Q hold15/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2821 VGND hold15/a_285_47# hold15/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2822 hold15/X hold15/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2823 VGND _257_/Q hold15/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2824 VPWR hold15/a_285_47# hold15/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2825 hold15/a_285_47# hold15/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2826 hold15/a_285_47# hold15/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2827 hold15/X hold15/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2864 VPWR tt_um_mult_4_22/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2865 uio_out[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2868 _219_/a_226_47# _218_/Y _219_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X2869 _219_/a_489_413# hold17/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2870 _219_/a_226_297# _208_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X2871 VPWR _216_/B _219_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2872 _219_/a_489_413# _219_/a_226_47# _219_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2873 _219_/a_76_199# _219_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X2874 VGND hold17/X _219_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2875 _219_/a_556_47# _216_/B _219_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2876 VGND _218_/Y _219_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2877 _219_/a_226_47# _208_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2878 VPWR _219_/a_76_199# _280_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X2879 VGND _219_/a_76_199# _280_/D VGND sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2924 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2925 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2926 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2927 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2928 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2929 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2930 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2931 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2932 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2933 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2934 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2935 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2936 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2937 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2938 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2939 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2940 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2941 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2942 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2943 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2944 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2945 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X2946 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2947 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2948 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2949 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2950 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2951 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2952 VGND clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2953 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2954 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2955 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2956 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2957 VPWR clkbuf_0_clk/a_110_47# clkbuf_0_clk/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2958 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2959 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2960 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2961 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2962 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2963 clkbuf_0_clk/X clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3100 VGND _270_/Q _183_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3101 _183_/a_68_297# _269_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3102 _202_/B _183_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3103 VPWR _270_/Q _183_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3104 _202_/B _183_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3105 _183_/a_150_297# _269_/Q _183_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3166 _166_/a_240_47# uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X3167 _276_/D _166_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3168 VGND _178_/A _166_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3169 _166_/a_51_297# _165_/X _166_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X3170 _166_/a_149_47# _186_/A _166_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X3171 _166_/a_240_47# _164_/Y _166_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3172 VPWR _178_/A _166_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3173 _276_/D _166_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X3174 _166_/a_149_47# _165_/X _166_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3175 _166_/a_245_297# _164_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3176 VPWR _186_/A _166_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3177 _166_/a_512_297# uo_out[5] _166_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3198 VPWR _263_/Q hold16/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3199 VGND hold16/a_285_47# hold16/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3200 hold16/X hold16/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3201 VGND _263_/Q hold16/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3202 VPWR hold16/a_285_47# hold16/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3203 hold16/a_285_47# hold16/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3204 hold16/a_285_47# hold16/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3205 hold16/X hold16/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3248 VPWR tt_um_mult_4_23/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3249 uio_out[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3250 _218_/a_377_297# _279_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X3251 _218_/a_47_47# _280_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X3252 _218_/a_129_47# _280_/Q _218_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3253 _218_/a_285_47# _280_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3254 _218_/Y _218_/a_47_47# _218_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X3255 VGND _279_/Q _218_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X3256 VPWR _279_/Q _218_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X3257 VPWR _218_/a_47_47# _218_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X3258 _218_/Y _280_/Q _218_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X3259 _218_/a_285_47# _279_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3262 VPWR uo_out[3] _149_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3263 _149_/Y uo_out[3] _149_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3264 _149_/a_113_47# _257_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3265 _149_/Y _257_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3350 _255_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3351 VGND _285_/CLK _255_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3352 _255_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3353 VPWR _285_/CLK _255_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3380 VPWR clkbuf_0_clk/X clkbuf_2_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3381 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3382 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3383 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3384 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3385 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3386 clkbuf_2_0__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3387 clkbuf_2_0__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3388 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3389 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3390 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3391 clkbuf_2_0__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3392 VGND clkbuf_0_clk/X clkbuf_2_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3393 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3394 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3395 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3396 VGND clkbuf_0_clk/X clkbuf_2_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3397 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3398 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3399 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3400 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3401 clkbuf_2_0__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3402 VPWR clkbuf_0_clk/X clkbuf_2_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3403 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3404 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3405 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3406 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3407 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3408 VGND clkbuf_2_0__f_clk/a_110_47# _267_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3409 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3410 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3411 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3412 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3413 VPWR clkbuf_2_0__f_clk/a_110_47# _267_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3414 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3415 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3416 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3417 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3418 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3419 _267_/CLK clkbuf_2_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3460 _182_/Y _269_/Q _182_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3461 _182_/Y _269_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3462 _182_/a_27_297# _270_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3463 VGND _270_/Q _182_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3464 _182_/Y _270_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3465 VGND _269_/Q _182_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3466 VPWR _270_/Q _182_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3467 _182_/a_27_297# _269_/Q _182_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3520 _165_/a_465_47# _153_/A _165_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3521 VGND _153_/B _165_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3522 VPWR _151_/Y _165_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3523 _165_/a_297_297# _153_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3524 _165_/a_297_297# _153_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X3525 VPWR _155_/A _165_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3526 _165_/a_381_47# _155_/A _165_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X3527 _165_/a_297_297# _128_/Y _165_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3528 VPWR _165_/a_79_21# _165_/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3529 _165_/a_79_21# _128_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X3530 VGND _165_/a_79_21# _165_/X VGND sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X3531 _165_/a_561_47# _151_/Y _165_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3552 VPWR _280_/Q hold17/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3553 VGND hold17/a_285_47# hold17/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3554 hold17/X hold17/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3555 VGND _280_/Q hold17/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3556 VPWR hold17/a_285_47# hold17/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3557 hold17/a_285_47# hold17/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3558 hold17/a_285_47# hold17/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3559 hold17/X hold17/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3602 VPWR tt_um_mult_4_24/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3603 uio_out[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3604 _279_/D _208_/Y _217_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3605 VPWR _216_/Y _279_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3606 _217_/a_27_47# _208_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3607 _279_/D _216_/Y _217_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3608 _217_/a_109_297# _216_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3609 VGND _216_/A _217_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3612 VPWR _148_/A _148_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3613 VPWR _148_/C _148_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3614 _148_/a_181_47# _148_/B _148_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3615 VGND _148_/C _148_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3616 _148_/a_27_47# _148_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3617 _148_/X _148_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X3618 _148_/X _148_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3619 _148_/a_109_47# _148_/A _148_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3780 VGND _128_/Y _181_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X3781 _181_/a_510_47# _180_/X _181_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X3782 _181_/a_79_21# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X3783 VPWR _180_/X _181_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3784 _181_/a_79_21# _177_/A _181_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X3785 _181_/a_297_297# _128_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3786 _181_/a_79_21# _186_/A _181_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X3787 VPWR _181_/a_79_21# _271_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3788 VGND _181_/a_79_21# _271_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3789 _181_/a_215_47# _177_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3848 VPWR _230_/X _233_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X3849 _233_/a_297_47# _211_/A _233_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3850 _233_/a_297_47# _230_/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3851 VGND _232_/X _233_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X3852 VPWR _233_/a_79_21# _285_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X3853 _233_/a_79_21# _211_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X3854 _233_/a_382_297# _232_/X _233_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X3855 VGND _233_/a_79_21# _285_/D VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3856 _164_/Y _153_/B _164_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3857 _164_/Y _153_/B _164_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3858 VPWR _151_/Y _164_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3859 _164_/a_109_297# _153_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3860 _164_/a_381_47# _153_/A _164_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3861 _164_/a_109_297# _155_/A _164_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3862 _164_/a_109_47# _155_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3863 VGND _151_/Y _164_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
X3864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3888 VPWR _255_/Q hold18/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3889 VGND hold18/a_285_47# hold18/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3890 hold18/X hold18/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3891 VGND _255_/Q hold18/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3892 VPWR hold18/a_285_47# hold18/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X3893 hold18/a_285_47# hold18/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3894 hold18/a_285_47# hold18/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X3895 hold18/X hold18/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3936 VPWR tt_um_mult_4_25/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3937 uio_out[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3938 VPWR tt_um_mult_4_14/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3939 uio_oe[0] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3940 VPWR _216_/A _216_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3941 _216_/Y _216_/A _216_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3942 _216_/a_113_47# _216_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3943 _216_/Y _216_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3946 _148_/C _144_/Y _147_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X3947 VPWR _146_/A _148_/C VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X3948 _147_/a_27_47# _144_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X3949 _148_/C _146_/A _147_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3950 _147_/a_109_297# _177_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3951 VGND _177_/A _147_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4086 _263_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4087 VGND _285_/CLK _263_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4088 _263_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4089 VPWR _285_/CLK _263_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4136 _180_/a_81_21# uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4137 _180_/a_299_297# uo_out[0] _180_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4138 VPWR _180_/a_81_21# _180_/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4139 VPWR _268_/Q _180_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4140 VGND _180_/a_81_21# _180_/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4141 VGND _263_/Q _180_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4142 _180_/a_299_297# _263_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4143 _180_/a_384_47# _268_/Q _180_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4206 VPWR _301_/a_27_47# uio_out[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4207 uio_out[1] _301_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4208 VPWR _301_/A _301_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4209 uio_out[1] _301_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4210 VGND _301_/a_27_47# uio_out[1] VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4211 VGND _301_/A _301_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4216 VPWR _232_/B _232_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X4217 _232_/X _232_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X4218 _232_/a_297_47# _232_/a_27_413# _232_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X4219 _232_/X _232_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4220 _232_/a_207_413# _232_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X4221 VPWR _284_/Q _232_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X4222 VGND _232_/B _232_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X4223 _232_/a_27_413# _284_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4226 VGND _128_/Y _163_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4227 _163_/a_510_47# _162_/X _163_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4228 _163_/a_79_21# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4229 VPWR _162_/X _163_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4230 _163_/a_79_21# _161_/X _163_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4231 _163_/a_297_297# _128_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4232 _163_/a_79_21# _186_/A _163_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4233 VPWR _163_/a_79_21# _277_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4234 VGND _163_/a_79_21# _277_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4235 _163_/a_215_47# _161_/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4258 VPWR _256_/Q hold19/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4259 VGND hold19/a_285_47# hold19/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X4260 hold19/X hold19/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4261 VGND _256_/Q hold19/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4262 VPWR hold19/a_285_47# hold19/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X4263 hold19/a_285_47# hold19/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X4264 hold19/a_285_47# hold19/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X4265 hold19/X hold19/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4312 VPWR tt_um_mult_4_26/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4313 uio_out[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4314 VPWR tt_um_mult_4_15/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4315 uio_oe[1] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4316 _215_/a_226_47# _216_/B _215_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=1.26 w=0.42 l=0.15
X4317 _215_/a_489_413# _229_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X4318 _215_/a_226_297# _283_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4319 VPWR _270_/Q _215_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4320 _215_/a_489_413# _215_/a_226_47# _215_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4321 _215_/a_76_199# _215_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X4322 VGND _229_/A _215_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4323 _215_/a_556_47# _270_/Q _215_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4324 VGND _216_/B _215_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4325 _215_/a_226_47# _283_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4326 VPWR _215_/a_76_199# _270_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4327 VGND _215_/a_76_199# _270_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4330 VPWR _146_/A _177_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4331 _177_/B _146_/A _146_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4332 _146_/a_113_47# _146_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4333 _177_/B _146_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4488 VPWR fanout11/a_27_47# _186_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4489 _186_/A fanout11/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4490 VPWR _127_/Y fanout11/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4491 _186_/A fanout11/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X4492 VGND fanout11/a_27_47# _186_/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4493 VGND _127_/Y fanout11/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4548 VPWR _231_/a_505_21# _231_/a_535_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4549 _231_/a_505_21# _285_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4550 _231_/a_218_374# _285_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4551 VGND _231_/a_505_21# _231_/a_439_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4552 _231_/a_76_199# _231_/A0 _231_/a_218_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4553 _231_/a_505_21# _285_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4554 _231_/a_439_47# _231_/A0 _231_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4555 _231_/a_535_374# _264_/Q _231_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X4556 _231_/a_76_199# _264_/Q _231_/a_218_47# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4557 _231_/a_218_47# _285_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4558 VPWR _231_/a_76_199# _232_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4559 VGND _231_/a_76_199# _232_/B VGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4562 VGND _178_/A _162_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4563 _162_/a_68_297# uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4564 _162_/X _162_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4565 VPWR _178_/A _162_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4566 _162_/X _162_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4567 _162_/a_150_297# uo_out[6] _162_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4598 VPWR input1/a_75_212# _254_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4599 input1/a_75_212# rst_n VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4600 input1/a_75_212# rst_n VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4601 VGND input1/a_75_212# _254_/D VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4620 _214_/a_226_47# _213_/X _214_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=1.26 w=0.42 l=0.15
X4621 _214_/a_489_413# _229_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X4622 _214_/a_226_297# _254_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4623 VPWR _269_/Q _214_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4624 _214_/a_489_413# _214_/a_226_47# _214_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4625 _214_/a_76_199# _214_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X4626 VGND _229_/A _214_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4627 _214_/a_556_47# _269_/Q _214_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4628 VGND _213_/X _214_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4629 _214_/a_226_47# _254_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4630 VPWR _214_/a_76_199# _269_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4631 VGND _214_/a_76_199# _269_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4634 VPWR tt_um_mult_4_27/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4635 uio_out[6] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4636 VPWR tt_um_mult_4_16/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4637 uio_oe[2] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4642 VGND uo_out[1] _145_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4643 _145_/a_68_297# _255_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4644 _146_/B _145_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4645 VPWR uo_out[1] _145_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4646 _146_/B _145_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4647 _145_/a_150_297# _255_/Q _145_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4650 _258_/CLK _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4651 VGND _267_/CLK _258_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4652 _258_/CLK _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4653 VPWR _267_/CLK _258_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4688 _274_/CLK _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4689 VGND _267_/CLK _274_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4690 _274_/CLK _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4691 VPWR _267_/CLK _274_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4700 _128_/Y _178_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4701 VGND _178_/A _128_/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4702 _128_/Y _178_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4703 VPWR _178_/A _128_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4842 VPWR _127_/Y fanout12/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4843 VPWR fanout12/a_27_47# _203_/A1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4844 VGND _127_/Y fanout12/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X4845 _203_/A1 fanout12/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4846 _203_/A1 fanout12/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4847 VGND fanout12/a_27_47# _203_/A1 VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4912 _230_/a_109_93# _285_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4913 _230_/X _230_/a_209_311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X4914 _230_/a_109_93# _285_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4915 _230_/a_296_53# _230_/a_109_93# _230_/a_209_311# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X4916 VPWR _284_/Q _230_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X4917 _230_/a_368_53# _230_/B _230_/a_296_53# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4918 _230_/X _230_/a_209_311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X4919 _230_/a_209_311# _230_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X4920 VPWR _230_/a_109_93# _230_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X4921 VGND _284_/Q _230_/a_368_53# VGND sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X4922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4926 _161_/X _161_/a_35_297# _161_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X4927 _161_/X _161_/B _161_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X4928 _161_/a_35_297# _161_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4929 _161_/a_117_297# _161_/B _161_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4930 VPWR _161_/B _161_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4931 VGND _161_/A _161_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4932 VGND _161_/a_35_297# _161_/X VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X4933 _161_/a_285_297# _161_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4934 VPWR _161_/A _161_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4935 _161_/a_285_47# _161_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4974 VPWR input2/a_75_212# input2/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4975 input2/a_75_212# ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4976 input2/a_75_212# ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4977 VGND input2/a_75_212# input2/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4998 _213_/a_109_93# _284_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4999 _213_/a_215_53# _283_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5000 VGND _213_/a_109_93# _213_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5001 VGND _285_/Q _213_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X5002 VPWR _285_/Q _213_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5003 _213_/a_369_297# _283_/Q _213_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X5004 _213_/X _213_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X5005 _213_/a_297_297# _213_/a_109_93# _213_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X5006 _213_/a_109_93# _284_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5007 _213_/X _213_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X5008 VPWR tt_um_mult_4_28/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5009 uio_out[7] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5010 VPWR tt_um_mult_4_17/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5011 uio_oe[3] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5014 VPWR uo_out[1] _144_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5015 VGND uo_out[1] _144_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5016 _144_/a_109_297# _255_/Q _144_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5017 _144_/Y _255_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5068 _127_/Y _270_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5069 VGND _270_/Q _127_/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5070 _127_/Y _270_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5071 VPWR _270_/Q _127_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5186 VPWR fanout13/a_27_47# _178_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5187 _178_/A fanout13/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5188 VPWR _268_/Q fanout13/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5189 _178_/A fanout13/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X5190 VGND fanout13/a_27_47# _178_/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5191 VGND _268_/Q fanout13/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5262 _160_/a_240_47# _178_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5263 _278_/D _160_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5264 VGND uo_out[7] _160_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5265 _160_/a_51_297# _159_/X _160_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X5266 _160_/a_149_47# _186_/A _160_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X5267 _160_/a_240_47# _158_/Y _160_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5268 VPWR uo_out[7] _160_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5269 _278_/D _160_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X5270 _160_/a_149_47# _159_/X _160_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5271 _160_/a_245_297# _158_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5272 VPWR _186_/A _160_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5273 _160_/a_512_297# _178_/A _160_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5314 VPWR input3/a_75_212# input3/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5315 input3/a_75_212# ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5316 input3/a_75_212# ui_in[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5317 VGND input3/a_75_212# input3/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5342 VPWR _284_/D _212_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X5343 _212_/a_27_297# _229_/A _212_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X5344 VGND _284_/D _212_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X5345 _268_/D _212_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X5346 _212_/a_27_297# _229_/A _212_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5347 _212_/a_109_297# _284_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X5348 _212_/a_373_47# _284_/Q _212_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X5349 _268_/D _212_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X5350 _212_/a_109_297# hold10/X _212_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5351 _212_/a_109_47# hold10/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X5352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5354 VPWR tt_um_mult_4_18/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5355 uio_oe[4] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5356 VPWR uo_out[0] _177_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5357 _177_/A uo_out[0] _143_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5358 _143_/a_113_47# _263_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5359 _177_/A _263_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5608 VPWR input4/a_75_212# input4/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5609 input4/a_75_212# ui_in[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5610 input4/a_75_212# ui_in[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5611 VGND input4/a_75_212# input4/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5614 VPWR clkbuf_0_clk/X clkbuf_2_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5615 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5616 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5617 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5618 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5619 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5620 clkbuf_2_1__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5621 clkbuf_2_1__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5622 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5623 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5624 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5625 clkbuf_2_1__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5626 VGND clkbuf_0_clk/X clkbuf_2_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5627 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5628 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5629 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5630 VGND clkbuf_0_clk/X clkbuf_2_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5631 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5632 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5633 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5634 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5635 clkbuf_2_1__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5636 VPWR clkbuf_0_clk/X clkbuf_2_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5637 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5638 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5639 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5640 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5641 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5642 VGND clkbuf_2_1__f_clk/a_110_47# clkload1/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5643 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5644 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5645 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5646 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5647 VPWR clkbuf_2_1__f_clk/a_110_47# clkload1/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5648 clkload1/A clkbuf_2_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5649 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5650 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5651 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5652 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5653 clkload1/A clkbuf_2_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5676 VPWR _211_/A _211_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5677 VGND _211_/A _229_/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5678 _211_/a_109_297# _211_/B _229_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5679 _229_/A _211_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5682 VPWR tt_um_mult_4_19/HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5683 uio_oe[5] VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
X5684 VPWR uo_out[1] _146_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5685 _146_/A uo_out[1] _142_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5686 _142_/a_113_47# _255_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5687 _146_/A _255_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5942 VPWR input5/a_75_212# input5/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5943 input5/a_75_212# ui_in[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5944 input5/a_75_212# ui_in[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5945 VGND input5/a_75_212# input5/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5986 VPWR _211_/A _210_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5987 _284_/D _210_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5988 VGND _211_/A _210_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5989 _210_/a_59_75# _285_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5990 _284_/D _210_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5991 _210_/a_145_75# _285_/Q _210_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X5992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5996 VGND uo_out[2] _141_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5997 _141_/a_68_297# _256_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5998 _148_/B _141_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5999 VPWR uo_out[2] _141_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6000 _148_/B _141_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6001 _141_/a_150_297# _256_/Q _141_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6106 _266_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6107 VGND _285_/CLK _266_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6108 _266_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6109 VPWR _285_/CLK _266_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6248 VPWR input6/a_75_212# input6/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6249 input6/a_75_212# ui_in[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6250 input6/a_75_212# ui_in[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6251 VGND input6/a_75_212# input6/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6286 VPWR uo_out[2] _148_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6287 _148_/A uo_out[2] _140_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6288 _140_/a_113_47# _256_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6289 _148_/A _256_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6320 _269_/Q _269_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6321 _269_/a_891_413# _269_/a_193_47# _269_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6322 _269_/a_561_413# _269_/a_27_47# _269_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6323 VPWR _285_/CLK _269_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6324 _269_/Q _269_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6325 _269_/a_381_47# _269_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6326 VGND _269_/a_634_159# _269_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6327 VPWR _269_/a_891_413# _269_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6328 _269_/a_466_413# _269_/a_193_47# _269_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6329 VPWR _269_/a_634_159# _269_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6330 _269_/a_634_159# _269_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6331 _269_/a_634_159# _269_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6332 _269_/a_975_413# _269_/a_193_47# _269_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6333 VGND _269_/a_1059_315# _269_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6334 _269_/a_193_47# _269_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6335 _269_/a_891_413# _269_/a_27_47# _269_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6336 _269_/a_592_47# _269_/a_193_47# _269_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6337 VPWR _269_/a_1059_315# _269_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6338 _269_/a_1017_47# _269_/a_27_47# _269_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6339 _269_/a_193_47# _269_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6340 _269_/a_466_413# _269_/a_27_47# _269_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6341 VGND _269_/a_891_413# _269_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6342 _269_/a_381_47# _269_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6343 VGND _285_/CLK _269_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6556 _285_/Q _285_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6557 _285_/a_891_413# _285_/a_193_47# _285_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6558 _285_/a_561_413# _285_/a_27_47# _285_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6559 VPWR _285_/CLK _285_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6560 _285_/Q _285_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6561 _285_/a_381_47# _285_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6562 VGND _285_/a_634_159# _285_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6563 VPWR _285_/a_891_413# _285_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6564 _285_/a_466_413# _285_/a_193_47# _285_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6565 VPWR _285_/a_634_159# _285_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6566 _285_/a_634_159# _285_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6567 _285_/a_634_159# _285_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6568 _285_/a_975_413# _285_/a_193_47# _285_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6569 VGND _285_/a_1059_315# _285_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6570 _285_/a_193_47# _285_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6571 _285_/a_891_413# _285_/a_27_47# _285_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6572 _285_/a_592_47# _285_/a_193_47# _285_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6573 VPWR _285_/a_1059_315# _285_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6574 _285_/a_1017_47# _285_/a_27_47# _285_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6575 _285_/a_193_47# _285_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6576 _285_/a_466_413# _285_/a_27_47# _285_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6577 VGND _285_/a_891_413# _285_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6578 _285_/a_381_47# _285_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6579 VGND _285_/CLK _285_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6582 VPWR input7/a_75_212# input7/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6583 input7/a_75_212# ui_in[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6584 input7/a_75_212# ui_in[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6585 VGND input7/a_75_212# input7/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6652 _268_/Q _268_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6653 _268_/a_891_413# _268_/a_193_47# _268_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6654 _268_/a_561_413# _268_/a_27_47# _268_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6655 VPWR _284_/CLK _268_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6656 _268_/Q _268_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6657 _268_/a_381_47# _268_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6658 VGND _268_/a_634_159# _268_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6659 VPWR _268_/a_891_413# _268_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6660 _268_/a_466_413# _268_/a_193_47# _268_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6661 VPWR _268_/a_634_159# _268_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6662 _268_/a_634_159# _268_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6663 _268_/a_634_159# _268_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6664 _268_/a_975_413# _268_/a_193_47# _268_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6665 VGND _268_/a_1059_315# _268_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6666 _268_/a_193_47# _268_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6667 _268_/a_891_413# _268_/a_27_47# _268_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6668 _268_/a_592_47# _268_/a_193_47# _268_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6669 VPWR _268_/a_1059_315# _268_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6670 _268_/a_1017_47# _268_/a_27_47# _268_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6671 _268_/a_193_47# _268_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6672 _268_/a_466_413# _268_/a_27_47# _268_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6673 VGND _268_/a_891_413# _268_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6674 _268_/a_381_47# _268_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6675 VGND _284_/CLK _268_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6676 _199_/a_240_47# input5/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6677 _257_/D _199_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6678 VGND _203_/A1 _199_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6679 _199_/a_51_297# hold19/X _199_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6680 _199_/a_149_47# _198_/X _199_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6681 _199_/a_240_47# _186_/Y _199_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6682 VPWR _203_/A1 _199_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6683 _257_/D _199_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6684 _199_/a_149_47# hold19/X _199_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6685 _199_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6686 VPWR _198_/X _199_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6687 _199_/a_512_297# input5/X _199_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6736 VPWR input10/a_75_212# _231_/A0 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6737 input10/a_75_212# uio_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6738 input10/a_75_212# uio_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6739 VGND input10/a_75_212# _231_/A0 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6860 _254_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6861 VGND _285_/CLK _254_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6862 _254_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6863 VPWR _285_/CLK _254_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6930 _284_/Q _284_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6931 _284_/a_891_413# _284_/a_193_47# _284_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6932 _284_/a_561_413# _284_/a_27_47# _284_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6933 VPWR _284_/CLK _284_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6934 _284_/Q _284_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6935 _284_/a_381_47# _284_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6936 VGND _284_/a_634_159# _284_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6937 VPWR _284_/a_891_413# _284_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6938 _284_/a_466_413# _284_/a_193_47# _284_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6939 VPWR _284_/a_634_159# _284_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6940 _284_/a_634_159# _284_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6941 _284_/a_634_159# _284_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6942 _284_/a_975_413# _284_/a_193_47# _284_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6943 VGND _284_/a_1059_315# _284_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6944 _284_/a_193_47# _284_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6945 _284_/a_891_413# _284_/a_27_47# _284_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6946 _284_/a_592_47# _284_/a_193_47# _284_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6947 VPWR _284_/a_1059_315# _284_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6948 _284_/a_1017_47# _284_/a_27_47# _284_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6949 _284_/a_193_47# _284_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6950 _284_/a_466_413# _284_/a_27_47# _284_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6951 VGND _284_/a_891_413# _284_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6952 _284_/a_381_47# _284_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6953 VGND _284_/CLK _284_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6954 VPWR input8/a_75_212# input8/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6955 input8/a_75_212# ui_in[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6956 input8/a_75_212# ui_in[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6957 VGND input8/a_75_212# input8/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7008 _301_/A _267_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7009 _267_/a_891_413# _267_/a_193_47# _267_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7010 _267_/a_561_413# _267_/a_27_47# _267_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7011 VPWR _267_/CLK _267_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7012 _301_/A _267_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7013 _267_/a_381_47# _267_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7014 VGND _267_/a_634_159# _267_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7015 VPWR _267_/a_891_413# _267_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7016 _267_/a_466_413# _267_/a_193_47# _267_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7017 VPWR _267_/a_634_159# _267_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7018 _267_/a_634_159# _267_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7019 _267_/a_634_159# _267_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7020 _267_/a_975_413# _267_/a_193_47# _267_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7021 VGND _267_/a_1059_315# _267_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7022 _267_/a_193_47# _267_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7023 _267_/a_891_413# _267_/a_27_47# _267_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7024 _267_/a_592_47# _267_/a_193_47# _267_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7025 VPWR _267_/a_1059_315# _267_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7026 _267_/a_1017_47# _267_/a_27_47# _267_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7027 _267_/a_193_47# _267_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7028 _267_/a_466_413# _267_/a_27_47# _267_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7029 VGND _267_/a_891_413# _267_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7030 _267_/a_381_47# _267_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7031 VGND _267_/CLK _267_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7034 VGND _257_/Q _198_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7035 _198_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7036 _198_/X _198_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7037 VPWR _257_/Q _198_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7038 _198_/X _198_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7039 _198_/a_150_297# _202_/B _198_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7130 _276_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7131 VGND clkload1/A _276_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7132 _276_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7133 VPWR clkload1/A _276_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7260 _283_/Q _283_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7261 _283_/a_891_413# _283_/a_193_47# _283_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7262 _283_/a_561_413# _283_/a_27_47# _283_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7263 VPWR _284_/CLK _283_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7264 _283_/Q _283_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7265 _283_/a_381_47# _283_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7266 VGND _283_/a_634_159# _283_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7267 VPWR _283_/a_891_413# _283_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7268 _283_/a_466_413# _283_/a_193_47# _283_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7269 VPWR _283_/a_634_159# _283_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7270 _283_/a_634_159# _283_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7271 _283_/a_634_159# _283_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7272 _283_/a_975_413# _283_/a_193_47# _283_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7273 VGND _283_/a_1059_315# _283_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7274 _283_/a_193_47# _283_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7275 _283_/a_891_413# _283_/a_27_47# _283_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7276 _283_/a_592_47# _283_/a_193_47# _283_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7277 VPWR _283_/a_1059_315# _283_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7278 _283_/a_1017_47# _283_/a_27_47# _283_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7279 _283_/a_193_47# _283_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7280 _283_/a_466_413# _283_/a_27_47# _283_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7281 VGND _283_/a_891_413# _283_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7282 _283_/a_381_47# _283_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7283 VGND _284_/CLK _283_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7288 VPWR input9/a_75_212# input9/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X7289 input9/a_75_212# ui_in[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X7290 input9/a_75_212# ui_in[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X7291 VGND input9/a_75_212# input9/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X7292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7338 hold7/A _266_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7339 _266_/a_891_413# _266_/a_193_47# _266_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7340 _266_/a_561_413# _266_/a_27_47# _266_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7341 VPWR _266_/CLK _266_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7342 hold7/A _266_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7343 _266_/a_381_47# _266_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7344 VGND _266_/a_634_159# _266_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7345 VPWR _266_/a_891_413# _266_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7346 _266_/a_466_413# _266_/a_193_47# _266_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7347 VPWR _266_/a_634_159# _266_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7348 _266_/a_634_159# _266_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7349 _266_/a_634_159# _266_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7350 _266_/a_975_413# _266_/a_193_47# _266_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7351 VGND _266_/a_1059_315# _266_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7352 _266_/a_193_47# _266_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7353 _266_/a_891_413# _266_/a_27_47# _266_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7354 _266_/a_592_47# _266_/a_193_47# _266_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7355 VPWR _266_/a_1059_315# _266_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7356 _266_/a_1017_47# _266_/a_27_47# _266_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7357 _266_/a_193_47# _266_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7358 _266_/a_466_413# _266_/a_27_47# _266_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7359 VGND _266_/a_891_413# _266_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7360 _266_/a_381_47# _266_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7361 VGND _266_/CLK _266_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7362 VPWR _182_/Y _197_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7363 _197_/a_27_297# _185_/X _197_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7364 VGND _182_/Y _197_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7365 _258_/D _197_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7366 _197_/a_27_297# _185_/X _197_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7367 _197_/a_109_297# hold12/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7368 _197_/a_373_47# hold12/X _197_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7369 _258_/D _197_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7370 _197_/a_109_297# hold15/X _197_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7371 _197_/a_109_47# hold15/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7524 VPWR hold1/A hold1/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7525 VGND hold1/a_285_47# hold1/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7526 hold1/X hold1/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7527 VGND hold1/A hold1/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7528 VPWR hold1/a_285_47# hold1/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7529 hold1/a_285_47# hold1/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7530 hold1/a_285_47# hold1/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7531 hold1/X hold1/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7632 hold4/A _282_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7633 _282_/a_891_413# _282_/a_193_47# _282_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7634 _282_/a_561_413# _282_/a_27_47# _282_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7635 VPWR _284_/CLK _282_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7636 hold4/A _282_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7637 _282_/a_381_47# _282_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7638 VGND _282_/a_634_159# _282_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7639 VPWR _282_/a_891_413# _282_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7640 _282_/a_466_413# _282_/a_193_47# _282_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7641 VPWR _282_/a_634_159# _282_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7642 _282_/a_634_159# _282_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7643 _282_/a_634_159# _282_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7644 _282_/a_975_413# _282_/a_193_47# _282_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7645 VGND _282_/a_1059_315# _282_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7646 _282_/a_193_47# _282_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7647 _282_/a_891_413# _282_/a_27_47# _282_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7648 _282_/a_592_47# _282_/a_193_47# _282_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7649 VPWR _282_/a_1059_315# _282_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7650 _282_/a_1017_47# _282_/a_27_47# _282_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7651 _282_/a_193_47# _282_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7652 _282_/a_466_413# _282_/a_27_47# _282_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7653 VGND _282_/a_891_413# _282_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7654 _282_/a_381_47# _282_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7655 VGND _284_/CLK _282_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7708 _265_/Q _265_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7709 _265_/a_891_413# _265_/a_193_47# _265_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7710 _265_/a_561_413# _265_/a_27_47# _265_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7711 VPWR _265_/CLK _265_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7712 _265_/Q _265_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7713 _265_/a_381_47# _265_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7714 VGND _265_/a_634_159# _265_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7715 VPWR _265_/a_891_413# _265_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7716 _265_/a_466_413# _265_/a_193_47# _265_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7717 VPWR _265_/a_634_159# _265_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7718 _265_/a_634_159# _265_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7719 _265_/a_634_159# _265_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7720 _265_/a_975_413# _265_/a_193_47# _265_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7721 VGND _265_/a_1059_315# _265_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7722 _265_/a_193_47# _265_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7723 _265_/a_891_413# _265_/a_27_47# _265_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7724 _265_/a_592_47# _265_/a_193_47# _265_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7725 VPWR _265_/a_1059_315# _265_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7726 _265_/a_1017_47# _265_/a_27_47# _265_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7727 _265_/a_193_47# _265_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7728 _265_/a_466_413# _265_/a_27_47# _265_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7729 VGND _265_/a_891_413# _265_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7730 _265_/a_381_47# _265_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7731 VGND _265_/CLK _265_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7732 VPWR _182_/Y _196_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7733 _196_/a_27_297# _185_/X _196_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7734 VGND _182_/Y _196_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7735 _259_/D _196_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7736 _196_/a_27_297# _185_/X _196_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7737 _196_/a_109_297# hold8/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7738 _196_/a_373_47# hold8/X _196_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7739 _259_/D _196_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7740 _196_/a_109_297# hold12/X _196_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7741 _196_/a_109_47# hold12/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7800 VGND _128_/Y _179_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X7801 _179_/a_510_47# _178_/X _179_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X7802 _179_/a_79_21# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X7803 VPWR _178_/X _179_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7804 _179_/a_79_21# _177_/X _179_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X7805 _179_/a_297_297# _128_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7806 _179_/a_79_21# _186_/A _179_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7807 VPWR _179_/a_79_21# _272_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7808 VGND _179_/a_79_21# _272_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7809 _179_/a_215_47# _177_/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7838 VPWR clkbuf_0_clk/X clkbuf_2_2__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7839 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7840 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7841 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7842 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7843 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7844 clkbuf_2_2__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7845 clkbuf_2_2__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7846 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7847 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7848 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7849 clkbuf_2_2__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7850 VGND clkbuf_0_clk/X clkbuf_2_2__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7851 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7852 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7853 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7854 VGND clkbuf_0_clk/X clkbuf_2_2__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7855 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7856 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7857 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7858 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7859 clkbuf_2_2__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7860 VPWR clkbuf_0_clk/X clkbuf_2_2__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7861 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7862 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7863 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7864 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7865 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7866 VGND clkbuf_2_2__f_clk/a_110_47# _284_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7867 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7868 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7869 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7870 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7871 VPWR clkbuf_2_2__f_clk/a_110_47# _284_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7872 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7873 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7874 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7875 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7876 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7877 _284_/CLK clkbuf_2_2__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7946 VPWR hold2/A hold2/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7947 VGND hold2/a_285_47# hold2/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7948 hold2/X hold2/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7949 VGND hold2/A hold2/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7950 VPWR hold2/a_285_47# hold2/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7951 hold2/a_285_47# hold2/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7952 hold2/a_285_47# hold2/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7953 hold2/X hold2/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7958 _256_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7959 VGND _285_/CLK _256_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7960 _256_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7961 VPWR _285_/CLK _256_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8048 hold5/A _281_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8049 _281_/a_891_413# _281_/a_193_47# _281_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8050 _281_/a_561_413# _281_/a_27_47# _281_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8051 VPWR _284_/CLK _281_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8052 hold5/A _281_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8053 _281_/a_381_47# _281_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8054 VGND _281_/a_634_159# _281_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8055 VPWR _281_/a_891_413# _281_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8056 _281_/a_466_413# _281_/a_193_47# _281_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8057 VPWR _281_/a_634_159# _281_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8058 _281_/a_634_159# _281_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8059 _281_/a_634_159# _281_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8060 _281_/a_975_413# _281_/a_193_47# _281_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8061 VGND _281_/a_1059_315# _281_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8062 _281_/a_193_47# _281_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8063 _281_/a_891_413# _281_/a_27_47# _281_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8064 _281_/a_592_47# _281_/a_193_47# _281_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8065 VPWR _281_/a_1059_315# _281_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8066 _281_/a_1017_47# _281_/a_27_47# _281_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8067 _281_/a_193_47# _281_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8068 _281_/a_466_413# _281_/a_27_47# _281_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8069 VGND _281_/a_891_413# _281_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8070 _281_/a_381_47# _281_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8071 VGND _284_/CLK _281_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8138 _264_/Q _264_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8139 _264_/a_891_413# _264_/a_193_47# _264_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8140 _264_/a_561_413# _264_/a_27_47# _264_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8141 VPWR _264_/CLK _264_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8142 _264_/Q _264_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8143 _264_/a_381_47# _264_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8144 VGND _264_/a_634_159# _264_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8145 VPWR _264_/a_891_413# _264_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8146 _264_/a_466_413# _264_/a_193_47# _264_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8147 VPWR _264_/a_634_159# _264_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8148 _264_/a_634_159# _264_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8149 _264_/a_634_159# _264_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8150 _264_/a_975_413# _264_/a_193_47# _264_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8151 VGND _264_/a_1059_315# _264_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8152 _264_/a_193_47# _264_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8153 _264_/a_891_413# _264_/a_27_47# _264_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8154 _264_/a_592_47# _264_/a_193_47# _264_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8155 VPWR _264_/a_1059_315# _264_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8156 _264_/a_1017_47# _264_/a_27_47# _264_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8157 _264_/a_193_47# _264_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8158 _264_/a_466_413# _264_/a_27_47# _264_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8159 VGND _264_/a_891_413# _264_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8160 _264_/a_381_47# _264_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8161 VGND _264_/CLK _264_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8162 VPWR _182_/Y _195_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8163 _195_/a_27_297# _185_/X _195_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8164 VGND _182_/Y _195_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8165 hold9/A _195_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8166 _195_/a_27_297# _185_/X _195_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8167 _195_/a_109_297# _260_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8168 _195_/a_373_47# _260_/Q _195_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8169 hold9/A _195_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8170 _195_/a_109_297# hold8/X _195_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8171 _195_/a_109_47# hold8/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8210 _273_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8211 VGND clkload1/A _273_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8212 _273_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8213 VPWR clkload1/A _273_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8236 VGND _178_/A _178_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8237 _178_/a_68_297# uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8238 _178_/X _178_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8239 VPWR _178_/A _178_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8240 _178_/X _178_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8241 _178_/a_150_297# uo_out[1] _178_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8322 VPWR hold3/A hold3/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8323 VGND hold3/a_285_47# hold3/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8324 hold3/X hold3/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8325 VGND hold3/A hold3/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8326 VPWR hold3/a_285_47# hold3/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8327 hold3/a_285_47# hold3/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8328 hold3/a_285_47# hold3/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8329 hold3/X hold3/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8406 _280_/Q _280_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8407 _280_/a_891_413# _280_/a_193_47# _280_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8408 _280_/a_561_413# _280_/a_27_47# _280_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8409 VPWR _284_/CLK _280_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8410 _280_/Q _280_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8411 _280_/a_381_47# _280_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8412 VGND _280_/a_634_159# _280_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8413 VPWR _280_/a_891_413# _280_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8414 _280_/a_466_413# _280_/a_193_47# _280_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8415 VPWR _280_/a_634_159# _280_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8416 _280_/a_634_159# _280_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8417 _280_/a_634_159# _280_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8418 _280_/a_975_413# _280_/a_193_47# _280_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8419 VGND _280_/a_1059_315# _280_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8420 _280_/a_193_47# _280_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8421 _280_/a_891_413# _280_/a_27_47# _280_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8422 _280_/a_592_47# _280_/a_193_47# _280_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8423 VPWR _280_/a_1059_315# _280_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8424 _280_/a_1017_47# _280_/a_27_47# _280_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8425 _280_/a_193_47# _280_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8426 _280_/a_466_413# _280_/a_27_47# _280_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8427 VGND _280_/a_891_413# _280_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8428 _280_/a_381_47# _280_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8429 VGND _284_/CLK _280_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8482 _263_/Q _263_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8483 _263_/a_891_413# _263_/a_193_47# _263_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8484 _263_/a_561_413# _263_/a_27_47# _263_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8485 VPWR _263_/CLK _263_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8486 _263_/Q _263_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8487 _263_/a_381_47# _263_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8488 VGND _263_/a_634_159# _263_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8489 VPWR _263_/a_891_413# _263_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8490 _263_/a_466_413# _263_/a_193_47# _263_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8491 VPWR _263_/a_634_159# _263_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8492 _263_/a_634_159# _263_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8493 _263_/a_634_159# _263_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8494 _263_/a_975_413# _263_/a_193_47# _263_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8495 VGND _263_/a_1059_315# _263_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8496 _263_/a_193_47# _263_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8497 _263_/a_891_413# _263_/a_27_47# _263_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8498 _263_/a_592_47# _263_/a_193_47# _263_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8499 VPWR _263_/a_1059_315# _263_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8500 _263_/a_1017_47# _263_/a_27_47# _263_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8501 _263_/a_193_47# _263_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8502 _263_/a_466_413# _263_/a_27_47# _263_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8503 VGND _263_/a_891_413# _263_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8504 _263_/a_381_47# _263_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8505 VGND _263_/CLK _263_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8508 VPWR _182_/Y _194_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8509 _194_/a_27_297# _185_/X _194_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8510 VGND _182_/Y _194_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8511 hold3/A _194_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8512 _194_/a_27_297# _185_/X _194_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8513 _194_/a_109_297# hold2/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8514 _194_/a_373_47# hold2/X _194_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8515 hold3/A _194_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8516 _194_/a_109_297# _260_/Q _194_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8517 _194_/a_109_47# _260_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8572 _177_/X _177_/a_35_297# _177_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8573 _177_/X _177_/B _177_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8574 _177_/a_35_297# _177_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8575 _177_/a_117_297# _177_/B _177_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8576 VPWR _177_/B _177_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8577 VGND _177_/A _177_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8578 VGND _177_/a_35_297# _177_/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8579 _177_/a_285_297# _177_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8580 VPWR _177_/A _177_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8581 _177_/a_285_47# _177_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8632 VPWR _229_/A _229_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8633 VGND _229_/A _283_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8634 _229_/a_109_297# _229_/B _283_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8635 _283_/D _229_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8676 VPWR hold4/A hold4/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8677 VGND hold4/a_285_47# hold4/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8678 hold4/X hold4/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8679 VGND hold4/A hold4/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8680 VPWR hold4/a_285_47# hold4/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8681 hold4/a_285_47# hold4/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8682 hold4/a_285_47# hold4/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8683 hold4/X hold4/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8836 hold1/A _262_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8837 _262_/a_891_413# _262_/a_193_47# _262_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8838 _262_/a_561_413# _262_/a_27_47# _262_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8839 VPWR _262_/CLK _262_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8840 hold1/A _262_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8841 _262_/a_381_47# _262_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8842 VGND _262_/a_634_159# _262_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8843 VPWR _262_/a_891_413# _262_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8844 _262_/a_466_413# _262_/a_193_47# _262_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8845 VPWR _262_/a_634_159# _262_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8846 _262_/a_634_159# _262_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8847 _262_/a_634_159# _262_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8848 _262_/a_975_413# _262_/a_193_47# _262_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8849 VGND _262_/a_1059_315# _262_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8850 _262_/a_193_47# _262_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8851 _262_/a_891_413# _262_/a_27_47# _262_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8852 _262_/a_592_47# _262_/a_193_47# _262_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8853 VPWR _262_/a_1059_315# _262_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8854 _262_/a_1017_47# _262_/a_27_47# _262_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8855 _262_/a_193_47# _262_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8856 _262_/a_466_413# _262_/a_27_47# _262_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8857 VGND _262_/a_891_413# _262_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8858 _262_/a_381_47# _262_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8859 VGND _262_/CLK _262_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8860 VPWR input9/X _193_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8861 _193_/a_27_297# _182_/Y _193_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8862 VGND input9/X _193_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8863 _262_/D _193_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8864 _193_/a_27_297# _182_/Y _193_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8865 _193_/a_109_297# _270_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8866 _193_/a_373_47# _270_/Q _193_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8867 _262_/D _193_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8868 _193_/a_109_297# hold1/X _193_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8869 _193_/a_109_47# hold1/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8934 VGND _178_/A _176_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8935 _176_/a_510_47# _175_/Y _176_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8936 _176_/a_79_21# _203_/A1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8937 VPWR _175_/Y _176_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8938 _176_/a_79_21# uo_out[2] _176_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8939 _176_/a_297_297# _178_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8940 _176_/a_79_21# _203_/A1 _176_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8941 VPWR _176_/a_79_21# _273_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8942 VGND _176_/a_79_21# _273_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8943 _176_/a_215_47# uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8958 _278_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8959 VGND clkload1/A _278_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8960 _278_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8961 VPWR clkload1/A _278_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9004 _228_/a_78_199# _227_/Y _228_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9005 VPWR _213_/X _228_/a_493_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X9006 _228_/a_493_297# _230_/B _228_/a_78_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X9007 VPWR _228_/a_78_199# _229_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X9008 VGND _230_/B _228_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X9009 _228_/a_78_199# _207_/X _228_/a_292_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X9010 _228_/a_215_47# _213_/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9011 _228_/a_215_47# _207_/X _228_/a_78_199# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X9012 _228_/a_292_297# _227_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9013 VGND _228_/a_78_199# _229_/B VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9016 _159_/a_81_21# _128_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X9017 _159_/a_299_297# _128_/Y _159_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X9018 VPWR _159_/a_81_21# _159_/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X9019 VPWR _158_/A _159_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9020 VGND _159_/a_81_21# _159_/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X9021 VGND _158_/B _159_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X9022 _159_/a_299_297# _158_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9023 _159_/a_384_47# _158_/A _159_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9068 VPWR hold5/A hold5/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9069 VGND hold5/a_285_47# hold5/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9070 hold5/X hold5/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9071 VGND hold5/A hold5/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9072 VPWR hold5/a_285_47# hold5/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9073 hold5/a_285_47# hold5/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9074 hold5/a_285_47# hold5/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9075 hold5/X hold5/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9208 hold2/A _261_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9209 _261_/a_891_413# _261_/a_193_47# _261_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X9210 _261_/a_561_413# _261_/a_27_47# _261_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X9211 VPWR _261_/CLK _261_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X9212 hold2/A _261_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9213 _261_/a_381_47# hold3/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X9214 VGND _261_/a_634_159# _261_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X9215 VPWR _261_/a_891_413# _261_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X9216 _261_/a_466_413# _261_/a_193_47# _261_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9217 VPWR _261_/a_634_159# _261_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9218 _261_/a_634_159# _261_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X9219 _261_/a_634_159# _261_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X9220 _261_/a_975_413# _261_/a_193_47# _261_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X9221 VGND _261_/a_1059_315# _261_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X9222 _261_/a_193_47# _261_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X9223 _261_/a_891_413# _261_/a_27_47# _261_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9224 _261_/a_592_47# _261_/a_193_47# _261_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X9225 VPWR _261_/a_1059_315# _261_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9226 _261_/a_1017_47# _261_/a_27_47# _261_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X9227 _261_/a_193_47# _261_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X9228 _261_/a_466_413# _261_/a_27_47# _261_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X9229 VGND _261_/a_891_413# _261_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X9230 _261_/a_381_47# hold3/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9231 VGND _261_/CLK _261_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9232 VPWR input2/X _192_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X9233 _192_/a_27_297# _182_/Y _192_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X9234 VGND input2/X _192_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X9235 _263_/D _192_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9236 _192_/a_27_297# _182_/Y _192_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X9237 _192_/a_109_297# _270_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9238 _192_/a_373_47# _270_/Q _192_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9239 _263_/D _192_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9240 _192_/a_109_297# hold16/X _192_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9241 _192_/a_109_47# hold16/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9296 _175_/Y _174_/Y _175_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X9297 VPWR _178_/A _175_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X9298 _175_/a_27_47# _174_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X9299 _175_/Y _178_/A _175_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9300 _175_/a_109_297# _148_/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9301 VGND _148_/X _175_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9310 _259_/CLK _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X9311 VGND _267_/CLK _259_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X9312 _259_/CLK _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9313 VPWR _267_/CLK _259_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9352 _227_/a_199_47# _218_/Y _227_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X9353 _227_/a_113_297# _222_/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X9354 _227_/Y _224_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X9355 VPWR _218_/Y _227_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X9356 _227_/a_113_297# _224_/Y _227_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9357 VGND _222_/X _227_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
X9358 VPWR _158_/A _158_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X9359 VGND _158_/A _158_/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X9360 _158_/a_109_297# _158_/B _158_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X9361 _158_/Y _158_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9396 VPWR hold7/A hold6/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9397 VGND hold6/a_285_47# hold6/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9398 hold6/X hold6/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9399 VGND hold7/A hold6/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9400 VPWR hold6/a_285_47# hold6/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9401 hold6/a_285_47# hold6/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9402 hold6/a_285_47# hold6/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9403 hold6/X hold6/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9532 _260_/Q _260_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9533 _260_/a_891_413# _260_/a_193_47# _260_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X9534 _260_/a_561_413# _260_/a_27_47# _260_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X9535 VPWR _260_/CLK _260_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X9536 _260_/Q _260_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9537 _260_/a_381_47# hold9/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X9538 VGND _260_/a_634_159# _260_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X9539 VPWR _260_/a_891_413# _260_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X9540 _260_/a_466_413# _260_/a_193_47# _260_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9541 VPWR _260_/a_634_159# _260_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9542 _260_/a_634_159# _260_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X9543 _260_/a_634_159# _260_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X9544 _260_/a_975_413# _260_/a_193_47# _260_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X9545 VGND _260_/a_1059_315# _260_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X9546 _260_/a_193_47# _260_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X9547 _260_/a_891_413# _260_/a_27_47# _260_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9548 _260_/a_592_47# _260_/a_193_47# _260_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X9549 VPWR _260_/a_1059_315# _260_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9550 _260_/a_1017_47# _260_/a_27_47# _260_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X9551 _260_/a_193_47# _260_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X9552 _260_/a_466_413# _260_/a_27_47# _260_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X9553 VGND _260_/a_891_413# _260_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X9554 _260_/a_381_47# hold9/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9555 VGND _260_/CLK _260_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9556 _191_/a_240_47# input6/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X9557 _264_/D _191_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X9558 VGND _203_/A1 _191_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9559 _191_/a_51_297# hold11/X _191_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X9560 _191_/a_149_47# _190_/X _191_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X9561 _191_/a_240_47# _186_/Y _191_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9562 VPWR _203_/A1 _191_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X9563 _264_/D _191_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X9564 _191_/a_149_47# hold11/X _191_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9565 _191_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9566 VPWR _190_/X _191_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9567 _191_/a_512_297# input6/X _191_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9624 _174_/a_199_47# _148_/A _174_/Y VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X9625 _174_/a_113_297# _148_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X9626 _174_/Y _148_/C VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9627 VPWR _148_/A _174_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9628 _174_/a_113_297# _148_/C _174_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X9629 VGND _148_/B _174_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9666 _265_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X9667 VGND _285_/CLK _265_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X9668 _265_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9669 VPWR _285_/CLK _265_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9688 _226_/a_27_297# _265_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9689 _226_/a_27_297# hold1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9690 _226_/a_277_297# _265_/Q _226_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9691 VPWR hold7/A _226_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X9692 _230_/B _226_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X9693 _226_/a_205_297# _264_/Q _226_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X9694 _230_/B _226_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X9695 VGND _264_/Q _226_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X9696 _226_/a_109_297# hold1/A _226_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9697 VGND hold7/A _226_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X9698 _158_/B _157_/a_35_297# _157_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X9699 _158_/B hold2/A _157_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X9700 _157_/a_35_297# hold2/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X9701 _157_/a_117_297# hold2/A _157_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X9702 VPWR hold2/A _157_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9703 VGND uo_out[7] _157_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9704 VGND _157_/a_35_297# _158_/B VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9705 _157_/a_285_297# uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9706 VPWR uo_out[7] _157_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9707 _157_/a_285_47# uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9712 _261_/CLK _267_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X9713 VGND _267_/CLK _261_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X9714 _261_/CLK _267_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9715 VPWR _267_/CLK _261_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9744 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9746 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9747 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9750 VPWR hold7/A hold7/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9751 VGND hold7/a_285_47# hold7/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9752 hold7/X hold7/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X9753 VGND hold7/A hold7/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9754 VPWR hold7/a_285_47# hold7/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X9755 hold7/a_285_47# hold7/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9756 hold7/a_285_47# hold7/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X9757 hold7/X hold7/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9774 _209_/a_222_93# _211_/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X9775 VPWR hold13/X _209_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9776 VGND _209_/a_79_199# _267_/D VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X9777 _209_/a_222_93# _211_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X9778 VGND _211_/B _209_/a_448_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X9779 _209_/a_448_47# _209_/a_222_93# _209_/a_79_199# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X9780 _209_/a_79_199# _209_/a_222_93# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X9781 _209_/a_544_297# _211_/B _209_/a_79_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X9782 _209_/a_448_47# hold13/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9783 VPWR _209_/a_79_199# _267_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X9784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9908 VGND _264_/Q _190_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X9909 _190_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X9910 _190_/X _190_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X9911 VPWR _264_/Q _190_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X9912 _190_/X _190_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X9913 _190_/a_150_297# _202_/B _190_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X9914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9978 VGND _178_/A _173_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X9979 _173_/a_510_47# _172_/Y _173_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X9980 _173_/a_79_21# _186_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X9981 VPWR _172_/Y _173_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9982 _173_/a_79_21# uo_out[3] _173_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X9983 _173_/a_297_297# _178_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X9984 _173_/a_79_21# _186_/A _173_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X9985 VPWR _173_/a_79_21# _274_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X9986 VGND _173_/a_79_21# _274_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X9987 _173_/a_215_47# uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X9988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X9991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X9992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X9993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X9994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X9995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X9996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X9998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X9999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10040 _225_/a_226_47# _208_/Y _225_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=1.26 w=0.42 l=0.15
X10041 _225_/a_489_413# _216_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X10042 _225_/a_226_297# _224_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10043 VPWR hold4/X _225_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10044 _225_/a_489_413# _225_/a_226_47# _225_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10045 _225_/a_76_199# _225_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X10046 VGND _216_/B _225_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10047 _225_/a_556_47# hold4/X _225_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10048 VGND _208_/Y _225_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10049 _225_/a_226_47# _224_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10050 VPWR _225_/a_76_199# _282_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X10051 VGND _225_/a_76_199# _282_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X10052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10054 _158_/A _133_/B _156_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.11863 ps=1.015 w=0.65 l=0.15
X10055 _156_/a_181_47# _155_/A _156_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X10056 VGND _131_/Y _158_/A VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10563 ps=0.975 w=0.65 l=0.15
X10057 VPWR _155_/A _156_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X10058 _158_/A _131_/Y _156_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X10059 _156_/a_109_297# _133_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X10060 _156_/a_109_297# _155_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10061 _156_/a_109_47# _155_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X10062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10104 VPWR hold8/A hold8/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10105 VGND hold8/a_285_47# hold8/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X10106 hold8/X hold8/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X10107 VGND hold8/A hold8/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10108 VPWR hold8/a_285_47# hold8/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X10109 hold8/a_285_47# hold8/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X10110 hold8/a_285_47# hold8/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X10111 hold8/X hold8/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X10112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10132 VPWR _283_/Q _208_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X10133 _208_/Y _283_/Q _208_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X10134 _208_/a_113_47# _211_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X10135 _208_/Y _211_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10140 VPWR _256_/Q _139_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10141 _139_/X _139_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X10142 VGND _256_/Q _139_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10143 _139_/a_59_75# uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10144 _139_/X _139_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X10145 _139_/a_145_75# uo_out[2] _139_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X10146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10190 VPWR clkbuf_0_clk/X clkbuf_2_3__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X10191 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X10192 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10193 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10194 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10195 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10196 clkbuf_2_3__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10197 clkbuf_2_3__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X10198 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X10199 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10200 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10201 clkbuf_2_3__f_clk/a_110_47# clkbuf_0_clk/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10202 VGND clkbuf_0_clk/X clkbuf_2_3__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10203 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10204 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10205 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10206 VGND clkbuf_0_clk/X clkbuf_2_3__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10207 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10208 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10209 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10210 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10211 clkbuf_2_3__f_clk/a_110_47# clkbuf_0_clk/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10212 VPWR clkbuf_0_clk/X clkbuf_2_3__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10213 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10214 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10215 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10216 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10217 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10218 VGND clkbuf_2_3__f_clk/a_110_47# _285_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10219 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10220 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10221 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10222 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10223 VPWR clkbuf_2_3__f_clk/a_110_47# _285_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10224 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10225 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10226 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10227 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10228 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10229 _285_/CLK clkbuf_2_3__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10334 VPWR _172_/B _172_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X10335 _172_/Y _178_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X10336 _172_/a_193_47# _172_/B _172_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X10337 _172_/Y _178_/A _172_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X10338 _172_/Y _172_/C VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10339 _172_/a_109_47# _172_/C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10360 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10361 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10384 _224_/a_377_297# hold4/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X10385 _224_/a_47_47# _224_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X10386 _224_/a_129_47# _224_/B _224_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X10387 _224_/a_285_47# _224_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X10388 _224_/Y _224_/a_47_47# _224_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X10389 VGND hold4/A _224_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X10390 VPWR hold4/A _224_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10391 VPWR _224_/a_47_47# _224_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X10392 _224_/Y _224_/B _224_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10393 _224_/a_285_47# hold4/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X10394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10398 VPWR _155_/A _161_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X10399 _161_/B _155_/A _155_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X10400 _155_/a_113_47# _155_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X10401 _161_/B _155_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10448 VPWR hold9/A hold9/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10449 VGND hold9/a_285_47# hold9/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X10450 hold9/X hold9/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X10451 VGND hold9/A hold9/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10452 VPWR hold9/a_285_47# hold9/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X10453 hold9/a_285_47# hold9/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X10454 hold9/a_285_47# hold9/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X10455 hold9/X hold9/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X10456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10464 _207_/a_109_93# _283_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X10465 _207_/a_215_53# _285_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X10466 VGND _207_/a_109_93# _207_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10467 VGND _284_/Q _207_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10468 VPWR _284_/Q _207_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1365 ps=1.49 w=0.42 l=0.15
X10469 _207_/a_369_297# _285_/Q _207_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X10470 _207_/X _207_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0 ps=0 w=1 l=0.15
X10471 _207_/a_297_297# _207_/a_109_93# _207_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10472 _207_/a_109_93# _283_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X10473 _207_/X _207_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X10474 VGND uo_out[3] _138_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10475 _138_/a_68_297# _257_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10476 _171_/B _138_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X10477 VPWR uo_out[3] _138_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X10478 _171_/B _138_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X10479 _138_/a_150_297# _257_/Q _138_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X10623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X10624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X10659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X10660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10668 VGND _151_/C _171_/a_27_93# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X10669 _172_/C _171_/a_27_93# _171_/a_206_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10670 _171_/a_206_47# _171_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X10671 VPWR _171_/a_27_93# _172_/C VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X10672 _172_/C _171_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X10673 VPWR _151_/C _171_/a_27_93# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X10674 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10678 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10679 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10683 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10685 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X10699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X10700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10722 _223_/a_226_47# _222_/X _223_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=1.26 w=0.42 l=0.15
X10723 _223_/a_489_413# hold5/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X10724 _223_/a_226_297# _208_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10725 VPWR _216_/B _223_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10726 _223_/a_489_413# _223_/a_226_47# _223_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X10727 _223_/a_76_199# _223_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X10728 VGND hold5/X _223_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10729 _223_/a_556_47# _216_/B _223_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10730 VGND _222_/X _223_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10731 _223_/a_226_47# _208_/Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10732 VPWR _223_/a_76_199# _281_/D VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X10733 VGND _223_/a_76_199# _281_/D VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X10734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10738 VPWR _154_/a_80_21# _155_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X10739 _154_/a_209_297# _151_/C VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X10740 _154_/a_303_47# _171_/B _154_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X10741 _154_/a_209_47# _151_/C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X10742 VGND _154_/a_80_21# _155_/B VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X10743 VGND _153_/Y _154_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X10744 _154_/a_80_21# _151_/A _154_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X10745 VPWR _171_/B _154_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X10746 _154_/a_80_21# _153_/Y _154_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X10747 _154_/a_209_297# _151_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X10748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10752 _275_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X10753 VGND clkload1/A _275_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X10754 _275_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X10755 VPWR clkload1/A _275_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X10756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10798 _216_/B _206_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X10799 _206_/a_111_297# _285_/Q _206_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X10800 _216_/B _206_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X10801 _206_/a_183_297# _284_/Q _206_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X10802 VPWR _254_/Q _206_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X10803 _206_/a_29_53# _284_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10804 VGND _285_/Q _206_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10805 VGND _254_/Q _206_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X10806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10808 VPWR _137_/B _137_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10809 _151_/A _137_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X10810 VGND _137_/B _137_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X10811 _137_/a_59_75# _153_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X10812 _151_/A _137_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X10813 _137_/a_145_75# _153_/A _137_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X10814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X10903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X10904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X10939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X10940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X10988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10990 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10996 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X10997 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X10998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X10999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11002 _170_/a_226_47# _148_/X _170_/a_226_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=1.26 w=0.42 l=0.15
X11003 _170_/a_489_413# _149_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X11004 _170_/a_226_297# _139_/X VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11005 VPWR _171_/B _170_/a_489_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11006 _170_/a_489_413# _170_/a_226_47# _170_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X11007 _170_/a_76_199# _170_/a_226_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X11008 VGND _149_/Y _170_/a_556_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X11009 _170_/a_556_47# _171_/B _170_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11010 VGND _148_/X _170_/a_226_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X11011 _170_/a_226_47# _139_/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11012 VPWR _170_/a_76_199# _172_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X11013 VGND _170_/a_76_199# _172_/B VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X11014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11034 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11035 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11036 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11037 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11048 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11049 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11050 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11051 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11057 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11066 VGND _224_/B _222_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X11067 _222_/a_68_297# _222_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11068 _222_/X _222_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X11069 VPWR _224_/B _222_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X11070 _222_/X _222_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X11071 _222_/a_150_297# _222_/B _222_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X11072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11080 VPWR _153_/A _153_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X11081 _153_/Y _153_/A _153_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X11082 _153_/a_113_47# _153_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11083 _153_/Y _153_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11088 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11089 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11090 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11103 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11134 VPWR _254_/Q _205_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11135 _205_/a_193_297# _284_/Q _205_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11136 _211_/B _284_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11137 VGND _254_/Q _211_/B VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X11138 _205_/a_109_297# _285_/Q _211_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11139 VGND _285_/Q _211_/B VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11144 VGND uo_out[4] _136_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X11145 _136_/a_68_297# _258_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11146 _137_/B _136_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X11147 VPWR uo_out[4] _136_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X11148 _137_/B _136_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X11149 _136_/a_150_297# _258_/Q _136_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X11150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11352 _221_/a_199_47# _279_/Q _222_/B VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X11353 _221_/a_113_297# _280_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X11354 _222_/B hold5/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11355 VPWR _279_/Q _221_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11356 _221_/a_113_297# hold5/A _222_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X11357 VGND _280_/Q _221_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11358 VPWR uo_out[5] _153_/B VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X11359 _153_/B uo_out[5] _152_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X11360 _152_/a_113_47# hold8/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11361 _153_/B hold8/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11364 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11366 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11373 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11375 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11379 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11380 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11381 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11398 VPWR _254_/Q _204_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X11399 VGND _254_/Q _211_/A VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X11400 _204_/a_109_297# _283_/Q _211_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X11401 _211_/A _283_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11404 VPWR uo_out[4] _153_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X11405 _153_/A uo_out[4] _135_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X11406 _135_/a_113_47# _258_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11407 _153_/A _258_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11424 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11425 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11429 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11432 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11433 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11434 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11435 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11514 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X11575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X11576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11618 _272_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X11619 VGND clkload1/A _272_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X11620 _272_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11621 VPWR clkload1/A _272_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11632 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11633 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11636 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11637 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11638 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11654 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11655 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11666 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11671 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11672 VPWR _279_/Q _220_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X11673 VPWR hold5/A _220_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11674 _220_/a_181_47# _280_/Q _220_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X11675 VGND hold5/A _220_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11676 _220_/a_27_47# _280_/Q VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11677 _224_/B _220_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X11678 _224_/B _220_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X11679 _220_/a_109_47# _279_/Q _220_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X11680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11682 VPWR _171_/B _151_/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X11683 _151_/Y _151_/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11684 _151_/a_193_47# _171_/B _151_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X11685 _151_/Y _151_/A _151_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X11686 _151_/Y _151_/C VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11687 _151_/a_109_47# _151_/C VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11699 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11700 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11708 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11709 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11718 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11719 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11720 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11721 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11726 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11728 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11729 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11730 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11740 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11742 _203_/a_240_47# input3/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X11743 _255_/D _203_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X11744 VGND _203_/A1 _203_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11745 _203_/a_51_297# hold20/X _203_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X11746 _203_/a_149_47# _202_/X _203_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X11747 _203_/a_240_47# _186_/Y _203_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11748 VPWR _203_/A1 _203_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X11749 _255_/D _203_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X11750 _203_/a_149_47# hold20/X _203_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X11751 _203_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11752 VPWR _202_/X _203_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11753 _203_/a_512_297# input3/X _203_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X11754 VGND uo_out[5] _134_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X11755 _134_/a_68_297# hold8/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X11756 _155_/A _134_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X11757 VPWR uo_out[5] _134_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X11758 _155_/A _134_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X11759 _134_/a_150_297# hold8/A _134_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X11760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11763 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11768 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11769 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11770 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11779 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11780 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11781 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11782 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11784 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11785 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11786 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11787 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11788 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11789 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11793 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11795 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11802 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11803 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11805 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11812 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11813 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11824 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11835 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11836 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11837 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11852 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11853 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11858 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11859 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11865 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11866 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11867 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11870 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11871 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11872 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11873 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11878 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11879 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11885 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11886 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11887 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11895 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11896 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11897 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11898 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11904 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11905 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11909 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11911 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11916 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11917 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11918 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11920 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11921 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11922 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11923 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11924 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11927 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11928 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11929 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11936 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11937 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11942 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11943 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11954 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11955 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11957 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11958 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X11961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X11962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X11965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X11966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11978 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11984 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11985 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11986 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X11987 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X11988 _150_/a_465_47# uo_out[3] _150_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11989 _151_/C _150_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X11990 _150_/a_109_297# _148_/B _150_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11991 _150_/a_193_297# _148_/C _150_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11992 _151_/C _150_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10238 ps=0.965 w=0.65 l=0.15
X11993 _150_/a_205_47# _148_/C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X11994 VPWR _257_/Q _150_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X11995 _150_/a_193_297# uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X11996 _150_/a_27_47# _148_/B _150_/a_205_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X11997 _150_/a_109_297# _139_/X _150_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11998 VGND _139_/X _150_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11999 VGND _257_/Q _150_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10238 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X12000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12010 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12011 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12019 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12024 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12025 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12026 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12027 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12032 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12033 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12034 _279_/Q _279_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X12035 _279_/a_891_413# _279_/a_193_47# _279_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X12036 _279_/a_561_413# _279_/a_27_47# _279_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X12037 VPWR _284_/CLK _279_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X12038 _279_/Q _279_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X12039 _279_/a_381_47# _279_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X12040 VGND _279_/a_634_159# _279_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X12041 VPWR _279_/a_891_413# _279_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X12042 _279_/a_466_413# _279_/a_193_47# _279_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12043 VPWR _279_/a_634_159# _279_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12044 _279_/a_634_159# _279_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X12045 _279_/a_634_159# _279_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X12046 _279_/a_975_413# _279_/a_193_47# _279_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X12047 VGND _279_/a_1059_315# _279_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X12048 _279_/a_193_47# _279_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X12049 _279_/a_891_413# _279_/a_27_47# _279_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12050 _279_/a_592_47# _279_/a_193_47# _279_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X12051 VPWR _279_/a_1059_315# _279_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12052 _279_/a_1017_47# _279_/a_27_47# _279_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X12053 _279_/a_193_47# _279_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X12054 _279_/a_466_413# _279_/a_27_47# _279_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X12055 VGND _279_/a_891_413# _279_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X12056 _279_/a_381_47# _279_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12057 VGND _284_/CLK _279_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X12058 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12060 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12061 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12070 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12072 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12073 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12074 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12075 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12076 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12080 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12081 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12088 VGND _255_/Q _202_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X12089 _202_/a_68_297# _202_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12090 _202_/X _202_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X12091 VPWR _255_/Q _202_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X12092 _202_/X _202_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X12093 _202_/a_150_297# _202_/B _202_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X12094 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12095 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12100 VPWR _133_/A _161_/A VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X12101 _161_/A _133_/A _133_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X12102 _133_/a_113_47# _133_/B VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12103 _161_/A _133_/B VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12104 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12106 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12108 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12112 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12113 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12114 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12116 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12117 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12120 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12121 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12122 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12123 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12125 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12126 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12128 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12129 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12132 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12133 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12135 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12136 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12137 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12139 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12147 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12148 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12149 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12151 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12153 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12162 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12164 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12165 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12182 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12183 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12187 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12190 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12191 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12207 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12208 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12209 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12213 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12214 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12216 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12218 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12219 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12245 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12246 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12247 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12251 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12263 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12264 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12265 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12266 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12267 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12268 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12269 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12270 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12271 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12282 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12298 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12299 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12300 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12306 _277_/CLK clkload1/A VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X12307 VGND clkload1/A _277_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X12308 _277_/CLK clkload1/A VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12309 VPWR clkload1/A _277_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12320 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12326 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12327 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12328 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12329 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12330 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12331 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12335 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12336 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12337 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12338 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12339 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12344 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12345 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12346 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12350 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12352 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12353 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12354 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12360 uo_out[7] _278_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0 ps=0 w=1 l=0.15
X12361 _278_/a_1020_47# _278_/a_27_47# _278_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.132 pd=1.49 as=0.1314 ps=1.45 w=0.36 l=0.15
X12362 _278_/a_572_47# _278_/a_193_47# _278_/a_475_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1374 pd=1.52 as=0.1188 ps=1.38 w=0.36 l=0.15
X12363 VPWR _278_/a_1062_300# _278_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1827 ps=1.71 w=0.42 l=0.15
X12364 _278_/a_634_183# _278_/a_475_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1978 pd=1.99 as=0 ps=0 w=0.64 l=0.15
X12365 VPWR _278_/CLK _278_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X12366 _278_/a_381_47# _278_/D VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0 ps=0 w=0.42 l=0.15
X12367 _278_/a_475_413# _278_/a_27_47# _278_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.36 l=0.15
X12368 VGND _278_/a_1062_300# _278_/a_1020_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12369 VPWR _278_/a_634_183# _278_/a_568_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X12370 uo_out[7] _278_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X12371 _278_/a_568_413# _278_/a_27_47# _278_/a_475_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1323 ps=1.47 w=0.42 l=0.15
X12372 _278_/a_634_183# _278_/a_475_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X12373 _278_/a_975_413# _278_/a_193_47# _278_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X12374 _278_/a_193_47# _278_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X12375 _278_/a_891_413# _278_/a_27_47# _278_/a_634_183# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12376 uo_out[7] _278_/a_1062_300# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12377 VGND _278_/a_891_413# _278_/a_1062_300# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X12378 VPWR _278_/a_1062_300# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12379 VGND _278_/a_1062_300# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12380 uo_out[7] _278_/a_1062_300# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12381 _278_/a_193_47# _278_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X12382 VGND _278_/a_1062_300# uo_out[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12383 _278_/a_381_47# _278_/D VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12384 VPWR _278_/a_891_413# _278_/a_1062_300# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X12385 _278_/a_475_413# _278_/a_193_47# _278_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12386 _278_/a_891_413# _278_/a_193_47# _278_/a_634_183# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X12387 VGND _278_/a_634_183# _278_/a_572_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12388 VGND _278_/CLK _278_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X12389 VPWR _278_/a_1062_300# uo_out[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12397 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12398 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12399 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12400 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12401 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12402 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12403 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12418 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12422 _201_/a_240_47# input4/X VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X12423 _256_/D _201_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X12424 VGND _203_/A1 _201_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12425 _201_/a_51_297# hold18/X _201_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X12426 _201_/a_149_47# _200_/X _201_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X12427 _201_/a_240_47# _186_/Y _201_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12428 VPWR _203_/A1 _201_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X12429 _256_/D _201_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X12430 _201_/a_149_47# hold18/X _201_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12431 _201_/a_245_297# _186_/Y VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12432 VPWR _200_/X _201_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12433 _201_/a_512_297# input4/X _201_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12434 VGND uo_out[6] _132_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X12435 _132_/a_68_297# _260_/Q VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12436 _133_/B _132_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X12437 VPWR uo_out[6] _132_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X12438 _133_/B _132_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X12439 _132_/a_150_297# _260_/Q _132_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X12440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12441 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12444 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12446 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12447 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12457 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12464 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12465 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12467 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12468 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12469 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12502 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12503 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12504 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12506 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12507 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12510 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12511 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12512 _257_/CLK _285_/CLK VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X12513 VGND _285_/CLK _257_/CLK VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X12514 _257_/CLK _285_/CLK VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X12515 VPWR _285_/CLK _257_/CLK VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X12516 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12517 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12518 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12520 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12526 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12528 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12529 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12539 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12542 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12543 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12546 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12548 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12549 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12553 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12568 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12578 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12579 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12580 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12581 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12584 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12585 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12589 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12591 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12596 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12597 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12598 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12599 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X12603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X12604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12608 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X12609 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X12610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12611 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12616 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12617 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12618 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12619 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X12627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X12628 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12629 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X12630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X12631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
