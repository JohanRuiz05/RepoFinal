* NGSPICE file created from tt_um_mult_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__dfxtp_4 VGND VPWR VNB VPB Q D CLK
X0 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X1 a_1020_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X2 a_572_47# a_193_47# a_475_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3 VPWR a_1062_300# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X4 a_634_183# a_475_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X5 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_475_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X8 VGND a_1062_300# a_1020_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X9 VPWR a_634_183# a_568_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09262 ps=0.935 w=0.65 l=0.15
X11 a_568_413# a_27_47# a_475_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X12 a_634_183# a_475_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X13 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_183# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 Q a_1062_300# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10563 ps=0.975 w=0.65 l=0.15
X17 VGND a_891_413# a_1062_300# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 Q a_1062_300# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 VGND a_1062_300# Q VNB sky130_fd_pr__nfet_01v8 ad=0.09262 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 VPWR a_891_413# a_1062_300# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X25 a_475_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X26 a_891_413# a_193_47# a_634_183# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X27 VGND a_634_183# a_572_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X29 VPWR a_1062_300# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__or2_1 VPB VNB VGND VPWR X A B
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 VPB VNB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 VPB VNB VGND VPWR A Y B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 X A VPB VNB VGND VPWR
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 VPB VNB VGND VPWR B1 B2 A2 A1 X C1
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_8 VNB VPB VGND VPWR A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1375 ps=1.275 w=1 l=0.15
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_2 VPB VNB VGND VPWR Y A B
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_6 VPB VNB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 VNB VPB VGND VPWR X A1 A2 B1 C1
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 Q CLK D VPB VNB VPWR VGND
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X20 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VPB VNB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_12 VNB VPB VGND VPWR Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.515 pd=3.03 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.33475 pd=2.33 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND VPB VNB A2 A1 B1 X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VNB VPB VGND VPWR B1 A1_N A2_N X B2
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VNB VPB VGND VPWR A X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VPB VNB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 VPB VNB VGND VPWR B Y A
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VPB VNB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 B1 Y A1 VPB VNB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 VPB VNB VGND VPWR A1 A2 B1 X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 VPWR VGND VPB VNB B2 B1 Y A1 A2
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VPB VNB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 X A_N B VGND VPWR VPB VNB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VPB VNB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VPB VNB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B X C VGND VPWR VPB VNB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 VNB VPB VPWR VGND A X B
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR VPB VNB B C_N A X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 VPB VNB VGND VPWR A B Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 VPB VNB VGND VPWR B2 A2 A1 B1 X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND VPB VNB B D C A X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VNB VPB VGND VPWR B1_N A1 A2 X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 VGND VPWR VPB VNB A3 A2 A1 Y B1
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.11863 ps=1.015 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10563 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1625 ps=1.325 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.1525 ps=1.305 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 VPB VNB VGND VPWR A B Y C
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 VPB VNB VGND VPWR A_N B Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 VPB VNB X A3 A2 A1 B1 VGND VPWR
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 VPB VNB VGND VPWR C B A Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND VPB VNB A1 A2 X B1 B2 C1
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10238 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10238 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
.ends

.subckt tt_um_mult_4 VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7]
XFILLER_67_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_77_169 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_277_ VGND VPWR VGND VPWR uo_out[6] _277_/D _277_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_10_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_200_ VPWR VGND VGND VPWR _200_/X _256_/Q _202_/B sky130_fd_sc_hd__or2_1
XFILLER_70_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_131_ VPWR VGND VPWR VGND _131_/Y _133_/A sky130_fd_sc_hd__inv_2
XFILLER_7_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_71_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_243__11 VPWR VGND VPWR VGND _264_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_77_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_46_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_41_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_276_ VGND VPWR VGND VPWR uo_out[5] _276_/D _276_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_10_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_43_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_130_ VPWR VGND VGND VPWR uo_out[6] _133_/A _260_/Q sky130_fd_sc_hd__nand2_1
XFILLER_7_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_259_ hold8/A _259_/CLK _259_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold20 hold20/X _263_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_35_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_46_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_275_ VGND VPWR VGND VPWR uo_out[4] _275_/D _275_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_69_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_64_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_258_ _258_/Q _258_/CLK _258_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_189_ VPWR VGND VGND VPWR _186_/Y hold6/X input7/X _203_/A1 _265_/D _188_/X sky130_fd_sc_hd__o221a_1
XFILLER_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_59_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_39_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold10 hold10/X _268_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_72_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_274_ VGND VPWR VGND VPWR uo_out[3] _274_/D _274_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_69_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_239__7 VPWR VGND VPWR VGND _260_/CLK _267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_36_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_46_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_257_ _257_/Q _257_/CLK _257_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_188_ VPWR VGND VGND VPWR _188_/X _265_/Q _202_/B sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_63_Left_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_75_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_47_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xhold11 hold11/X _265_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_273_ VGND VPWR VGND VPWR uo_out[2] _273_/D _273_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_6_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_256_ _256_/Q _256_/CLK _256_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_187_ VPWR VGND VGND VPWR _186_/Y hold1/X input8/X _186_/A _266_/D _184_/X sky130_fd_sc_hd__o221a_1
X_241__9 VPWR VGND VPWR VGND _262_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_669 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 VGND VPWR VGND VPWR _267_/CLK clkload0/Y sky130_fd_sc_hd__clkinv_8
XFILLER_7_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 hold12/X _258_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_274 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_37_Right_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_58_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_272_ VGND VPWR VGND VPWR uo_out[1] _272_/D _272_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_6_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_255_ _255_/Q _255_/CLK _255_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_64 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_186_ VPWR VGND VGND VPWR _186_/Y _186_/A _269_/Q sky130_fd_sc_hd__nand2_2
XFILLER_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 VPWR VGND VPWR VGND clkload1/Y clkload1/A sky130_fd_sc_hd__inv_6
XFILLER_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_169_ VGND VPWR VGND VPWR _275_/D _178_/A uo_out[4] _168_/X _186_/A sky130_fd_sc_hd__o211a_1
XFILLER_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold13 hold13/X _301_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_20 uio_oe[6] tt_um_mult_4_20/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_57_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Left_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_271_ uo_out[0] _271_/CLK _271_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_2
XFILLER_6_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_254_ _254_/Q _254_/CLK _254_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_80_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_185_ VPWR VGND _185_/X _269_/Q _186_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_56_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 VGND VPWR VGND VPWR clkload2/Y _284_/CLK sky130_fd_sc_hd__inv_12
XFILLER_59_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ VPWR VGND VPWR VGND _167_/X _151_/Y _128_/Y _168_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_38_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold14 _216_/A _279_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_21 uio_oe[7] tt_um_mult_4_21/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_246__14 VPWR VGND VPWR VGND _271_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ _270_/Q _284_/CLK _270_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_184_ VPWR VGND VGND VPWR _184_/X hold7/X _202_/B sky130_fd_sc_hd__or2_1
XFILLER_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_167_ VPWR VGND VPWR VGND _151_/C _171_/B _151_/A _167_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 hold15/X _257_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_22 uio_out[0] tt_um_mult_4_22/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_219_ VGND VPWR VGND VPWR hold17/X _208_/Y _218_/Y _280_/D _216_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk VGND VPWR VGND VPWR clk clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Right_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_54_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_91 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_63_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_45_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_183_ VPWR VGND VGND VPWR _202_/B _270_/Q _269_/Q sky130_fd_sc_hd__or2_1
XFILLER_6_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_239 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_74_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_166_ VPWR VGND VGND VPWR _164_/Y _165_/X uo_out[5] _178_/A _276_/D _186_/A sky130_fd_sc_hd__o221a_1
XFILLER_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 hold16/X _263_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_23 uio_out[2] tt_um_mult_4_23/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_218_ VGND VPWR _280_/Q _218_/Y _279_/Q VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_7_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_149_ VPWR VGND VGND VPWR uo_out[3] _149_/Y _257_/Q sky130_fd_sc_hd__nand2_1
XFILLER_7_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_234__2 VPWR VGND VPWR VGND _255_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_clk VGND VPWR VGND VPWR clkbuf_0_clk/X _267_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_57 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_182_ VPWR VGND VGND VPWR _269_/Q _182_/Y _270_/Q sky130_fd_sc_hd__nor2_2
XFILLER_13_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_192 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_165_ VGND VPWR _151_/Y _153_/B _153_/A _165_/X _128_/Y _155_/A VPWR VGND sky130_fd_sc_hd__a41o_1
XFILLER_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 hold17/X _280_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xtt_um_mult_4_24 uio_out[3] tt_um_mult_4_24/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_217_ VGND VPWR _208_/Y _216_/Y _279_/D _216_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_148_ VGND VPWR _148_/X _148_/B _148_/A _148_/C VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_7_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_57_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_181_ VGND VPWR VGND VPWR _271_/D _128_/Y _177_/A _180_/X _186_/A sky130_fd_sc_hd__o211a_1
XFILLER_10_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_47_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_233_ VPWR VGND VGND VPWR _230_/X _232_/X _211_/A _285_/D sky130_fd_sc_hd__o21a_1
X_164_ VPWR VGND VPWR VGND _155_/A _153_/B _164_/Y _153_/A _151_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_6_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 hold18/X _255_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_288 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_25 uio_out[4] tt_um_mult_4_25/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xtt_um_mult_4_14 uio_oe[0] tt_um_mult_4_14/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_216_ VPWR VGND VGND VPWR _216_/A _216_/Y _216_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_147_ VGND VPWR _144_/Y _146_/A _148_/C _177_/A VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_95 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_10_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_242__10 VPWR VGND VPWR VGND _263_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_72_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ VPWR VGND VPWR VGND _263_/Q _268_/Q uo_out[0] _180_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ VPWR VGND uio_out[1] _301_/A VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_232_ _232_/X _284_/Q _232_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__and2b_1
XFILLER_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_163_ VGND VPWR VGND VPWR _277_/D _128_/Y _161_/X _162_/X _186_/A sky130_fd_sc_hd__o211a_1
XFILLER_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xhold19 hold19/X _256_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_29_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_71_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_74_201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_27_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_42_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_26 uio_out[5] tt_um_mult_4_26/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xtt_um_mult_4_15 uio_oe[1] tt_um_mult_4_15/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_215_ VGND VPWR VGND VPWR _229_/A _283_/Q _216_/B _270_/D _270_/Q sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_146_ VPWR VGND VGND VPWR _146_/A _177_/B _146_/B sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_2_Left_83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_69_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_326 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_35_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout11 VPWR VGND _186_/A _127_/Y VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_10_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_231_ VGND VPWR VPWR VGND _232_/B _264_/Q _285_/Q _231_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_162_ VPWR VGND VGND VPWR _162_/X _178_/A uo_out[6] sky130_fd_sc_hd__or2_1
XFILLER_10_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 VGND VPWR _254_/D rst_n VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_37_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_214_ VGND VPWR VGND VPWR _229_/A _254_/Q _213_/X _269_/D _269_/Q sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_27 uio_out[6] tt_um_mult_4_27/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xtt_um_mult_4_16 uio_oe[2] tt_um_mult_4_16/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_145_ VPWR VGND VGND VPWR _146_/B uo_out[1] _255_/Q sky130_fd_sc_hd__or2_1
XFILLER_19_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_237__5 VPWR VGND VPWR VGND _258_/CLK _267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_249__17 VPWR VGND VPWR VGND _274_/CLK _267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_128_ VPWR VGND VPWR VGND _128_/Y _178_/A sky130_fd_sc_hd__inv_2
XFILLER_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_35_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_73_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_54_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_143 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_72_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout12 VGND VPWR _127_/Y _203_/A1 VPWR VGND sky130_fd_sc_hd__clkbuf_2
XFILLER_10_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_230_ _285_/Q _230_/B _230_/X _284_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__and3b_1
XFILLER_23_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_161_ VGND VPWR VPWR VGND _161_/A _161_/X _161_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_77_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_65_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput2 VGND VPWR input2/X ui_in[0] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_68_266 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_213_ VGND VPWR VPWR VGND _283_/Q _284_/Q _285_/Q _213_/X sky130_fd_sc_hd__or3b_1
Xtt_um_mult_4_28 uio_out[7] tt_um_mult_4_28/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
Xtt_um_mult_4_17 uio_oe[3] tt_um_mult_4_17/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_144_ VPWR VGND VGND VPWR uo_out[1] _255_/Q _144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_127_ VPWR VGND VPWR VGND _127_/Y _270_/Q sky130_fd_sc_hd__inv_2
XFILLER_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_66_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_35_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout13 VPWR VGND _178_/A _268_/Q VPWR VGND sky130_fd_sc_hd__buf_2
XFILLER_54_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_26_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ VPWR VGND VGND VPWR _158_/Y _159_/X _178_/A uo_out[7] _278_/D _186_/A sky130_fd_sc_hd__o221a_1
XFILLER_24_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_68_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput3 VGND VPWR input3/X ui_in[1] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_55_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_212_ VPWR VGND VPWR VGND _229_/A _284_/Q _284_/D _268_/D hold10/X sky130_fd_sc_hd__a22o_1
XFILLER_42_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xtt_um_mult_4_18 uio_oe[4] tt_um_mult_4_18/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_143_ VPWR VGND VGND VPWR uo_out[0] _177_/A _263_/Q sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_54_Right_54 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_65_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_63_Right_63 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_80_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Right_72 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_40_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_43_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_140 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 VGND VPWR input4/X ui_in[2] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_36_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_clk VGND VPWR VGND VPWR clkbuf_0_clk/X clkload1/A sky130_fd_sc_hd__clkbuf_16
XFILLER_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_211_ VPWR VGND VGND VPWR _211_/A _211_/B _229_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xtt_um_mult_4_19 uio_oe[5] tt_um_mult_4_19/HI VPWR VGND VGND VPWR sky130_fd_sc_hd__conb_1
X_142_ VPWR VGND VGND VPWR uo_out[1] _146_/A _255_/Q sky130_fd_sc_hd__nand2_1
XFILLER_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_16_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_66_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_22_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Left_112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_1_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput5 VGND VPWR input5/X ui_in[3] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_49_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_210_ VPWR VGND _284_/D _211_/A _285_/Q VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_70_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_141_ VPWR VGND VGND VPWR _148_/B uo_out[2] _256_/Q sky130_fd_sc_hd__or2_1
XFILLER_7_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_34_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_331 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_29_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_245__13 VPWR VGND VPWR VGND _266_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_69_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 VGND VPWR input6/X ui_in[4] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_49_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_140_ VPWR VGND VGND VPWR uo_out[2] _148_/A _256_/Q sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Right_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_78_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Right_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_269_ _269_/Q _285_/CLK _269_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_41_Right_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_67_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_285_ _285_/Q _285_/CLK _285_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_49_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput7 VGND VPWR input7/X ui_in[5] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_49_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_268_ _268_/Q _284_/CLK _268_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_199_ VPWR VGND VGND VPWR _186_/Y hold19/X input5/X _203_/A1 _257_/D _198_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_15_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_78_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput10 VGND VPWR _231_/A0 uio_in[0] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_57_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_44_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_94 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_129__1 VPWR VGND VPWR VGND _254_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_284_ _284_/Q _284_/CLK _284_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
Xinput8 VGND VPWR input8/X ui_in[6] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_267_ _301_/A _267_/CLK _267_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_10_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_198_ VPWR VGND VGND VPWR _198_/X _257_/Q _202_/B sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_47_Left_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_75_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_68_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_251__19 VPWR VGND VPWR VGND _276_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_3_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_283_ _283_/Q _284_/CLK _283_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 VGND VPWR input9/X ui_in[7] VPWR VGND sky130_fd_sc_hd__clkbuf_1
XFILLER_64_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ hold7/A _266_/CLK _266_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_197_ VPWR VGND VPWR VGND _185_/X hold12/X _182_/Y _258_/D hold15/X sky130_fd_sc_hd__a22o_1
XFILLER_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_47_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_47_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 hold1/X hold1/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_50_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_71_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_50_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ hold4/A _284_/CLK _282_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_69_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_265_ _265_/Q _265_/CLK _265_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_196_ VPWR VGND VPWR VGND _185_/X hold8/X _182_/Y _259_/D hold12/X sky130_fd_sc_hd__a22o_1
XFILLER_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_247 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_179_ VGND VPWR VGND VPWR _272_/D _128_/Y _177_/X _178_/X _186_/A sky130_fd_sc_hd__o211a_1
XFILLER_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_65_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk VGND VPWR VGND VPWR clkbuf_0_clk/X _284_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold2 hold2/X hold2/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_235__3 VPWR VGND VPWR VGND _256_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_76_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_98 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_281_ hold5/A _284_/CLK _281_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_264_ _264_/Q _264_/CLK _264_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_195_ VPWR VGND VPWR VGND _185_/X _260_/Q _182_/Y hold9/A hold8/X sky130_fd_sc_hd__a22o_1
XFILLER_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_64_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Left_106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_43_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_51_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_248__16 VPWR VGND VPWR VGND _273_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_52_Left_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ VPWR VGND VGND VPWR _178_/X _178_/A uo_out[1] sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_70_Left_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold3 hold3/X hold3/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_76_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _280_/Q _284_/CLK _280_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_268 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_263_ _263_/Q _263_/CLK _263_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XFILLER_6_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_194_ VPWR VGND VPWR VGND _185_/X hold2/X _182_/Y hold3/A _260_/Q sky130_fd_sc_hd__a22o_1
XFILLER_6_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_177_ VGND VPWR VPWR VGND _177_/A _177_/X _177_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_229_ VPWR VGND VGND VPWR _229_/A _229_/B _283_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 hold4/X hold4/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_62_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_8_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_73_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_50_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_262_ hold1/A _262_/CLK _262_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_193_ VPWR VGND VPWR VGND _182_/Y _270_/Q input9/X _262_/D hold1/X sky130_fd_sc_hd__a22o_1
XFILLER_6_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_176_ VGND VPWR VGND VPWR _273_/D _178_/A uo_out[2] _175_/Y _203_/A1 sky130_fd_sc_hd__o211a_1
XFILLER_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_253__21 VPWR VGND VPWR VGND _278_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_56_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_70_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ VPWR VGND VGND VPWR _207_/X _230_/B _213_/X _227_/Y _229_/B sky130_fd_sc_hd__o22a_1
XFILLER_7_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ VPWR VGND VPWR VGND _158_/B _158_/A _128_/Y _159_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 hold5/X hold5/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_58_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_261_ hold2/A _261_/CLK hold3/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_192_ VPWR VGND VPWR VGND _182_/Y _270_/Q input2/X _263_/D hold16/X sky130_fd_sc_hd__a22o_1
XFILLER_6_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_74_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Left_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_175_ VGND VPWR _174_/Y _178_/A _175_/Y _148_/X VPWR VGND sky130_fd_sc_hd__o21ai_1
XFILLER_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_238__6 VPWR VGND VPWR VGND _259_/CLK _267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_59_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_30_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ VPWR VGND VPWR VGND _222_/X _218_/Y _224_/Y _227_/Y sky130_fd_sc_hd__a21oi_1
X_158_ VPWR VGND VGND VPWR _158_/A _158_/B _158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 hold6/X hold7/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_79_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_26_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_216 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_260_ _260_/Q _260_/CLK hold9/X VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
X_191_ VPWR VGND VGND VPWR _186_/Y hold11/X input6/X _203_/A1 _264_/D _190_/X sky130_fd_sc_hd__o221a_1
XFILLER_10_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_27_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_174_ VPWR VGND VPWR VGND _148_/B _148_/A _148_/C _174_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_244__12 VPWR VGND VPWR VGND _265_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_74_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_226_ VPWR VGND VPWR VGND _265_/Q hold1/A _264_/Q hold7/A _230_/B sky130_fd_sc_hd__or4_1
X_157_ VGND VPWR VPWR VGND uo_out[7] _158_/B hold2/A sky130_fd_sc_hd__xor2_1
XFILLER_7_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_240__8 VPWR VGND VPWR VGND _261_/CLK _267_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xhold7 hold7/X hold7/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_209_ VGND VPWR VGND VPWR _211_/A hold13/X _211_/B _267_/D sky130_fd_sc_hd__o21ba_1
XFILLER_7_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_100 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_22_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_67_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_75_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_31_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_41_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_190_ VPWR VGND VGND VPWR _190_/X _264_/Q _202_/B sky130_fd_sc_hd__or2_1
XFILLER_50_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_173_ VGND VPWR VGND VPWR _274_/D _178_/A uo_out[3] _172_/Y _186_/A sky130_fd_sc_hd__o211a_1
XFILLER_6_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_77_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_37_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_80_529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_225_ VGND VPWR VGND VPWR _216_/B _224_/Y _208_/Y _282_/D hold4/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_156_ VGND VPWR VPWR VGND _155_/B _155_/A _133_/B _158_/A _131_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_81 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_61_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 hold8/X hold8/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_75_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_74_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_208_ VPWR VGND VGND VPWR _283_/Q _208_/Y _211_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_139_ VPWR VGND _139_/X _256_/Q uo_out[2] VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk VGND VPWR VGND VPWR clkbuf_0_clk/X _285_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_49_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ VPWR VGND VGND VPWR _178_/A _172_/B _172_/Y _172_/C sky130_fd_sc_hd__nand3_1
XFILLER_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_42_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_224_ VGND VPWR _224_/B _224_/Y hold4/A VPWR VGND sky130_fd_sc_hd__xnor2_1
XFILLER_11_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_155_ VPWR VGND VGND VPWR _155_/A _161_/B _155_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 hold9/X hold9/A VPWR VGND VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_207_ VGND VPWR VPWR VGND _285_/Q _283_/Q _284_/Q _207_/X sky130_fd_sc_hd__or3b_1
X_138_ VPWR VGND VGND VPWR _171_/B uo_out[3] _257_/Q sky130_fd_sc_hd__or2_1
XFILLER_7_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_38_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_57_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_171_ VPWR VGND VGND VPWR _151_/C _171_/B _172_/C sky130_fd_sc_hd__nand2b_1
XFILLER_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_79_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_223_ VGND VPWR VGND VPWR hold5/X _208_/Y _222_/X _281_/D _216_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_154_ VPWR VGND _155_/B _151_/C _171_/B _151_/A _153_/Y VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_11_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_250__18 VPWR VGND VPWR VGND _275_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_34_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_206_ VPWR VGND VPWR VGND _284_/Q _285_/Q _254_/Q _216_/B sky130_fd_sc_hd__or3_1
XFILLER_11_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_137_ VPWR VGND _151_/A _137_/B _153_/A VPWR VGND sky130_fd_sc_hd__and2_1
XFILLER_66_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_228 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_72_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_97 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_39_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ VGND VPWR VGND VPWR _149_/Y _139_/X _148_/X _172_/B _171_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_68_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_222_ VPWR VGND VGND VPWR _222_/X _224_/B _222_/B sky130_fd_sc_hd__or2_1
XFILLER_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_153_ VPWR VGND VGND VPWR _153_/A _153_/Y _153_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_85 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_205_ VPWR VGND VGND VPWR _285_/Q _284_/Q _254_/Q _211_/B sky130_fd_sc_hd__nor3_1
XFILLER_11_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_136_ VPWR VGND VGND VPWR _137_/B uo_out[4] _258_/Q sky130_fd_sc_hd__or2_1
XFILLER_66_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_40_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_26_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_73_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_68_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_221_ VPWR VGND VPWR VGND _280_/Q _279_/Q hold5/A _222_/B sky130_fd_sc_hd__a21oi_1
X_152_ VPWR VGND VGND VPWR uo_out[5] _153_/B hold8/A sky130_fd_sc_hd__nand2_1
XFILLER_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_204_ VPWR VGND VGND VPWR _254_/Q _283_/Q _211_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_135_ VPWR VGND VGND VPWR uo_out[4] _153_/A _258_/Q sky130_fd_sc_hd__nand2_1
XFILLER_11_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_19_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_69_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_123 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_132 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_59_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_27_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_72_244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_51_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_247__15 VPWR VGND VPWR VGND _272_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_2_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_70_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ VGND VPWR _224_/B _280_/Q _279_/Q hold5/A VPWR VGND sky130_fd_sc_hd__and3_1
XFILLER_23_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ VPWR VGND VGND VPWR _151_/A _171_/B _151_/Y _151_/C sky130_fd_sc_hd__nand3_1
XFILLER_10_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ VPWR VGND VGND VPWR _186_/Y hold20/X input3/X _203_/A1 _255_/D _202_/X sky130_fd_sc_hd__o221a_1
X_134_ VPWR VGND VGND VPWR _155_/A uo_out[5] hold8/A sky130_fd_sc_hd__or2_1
XFILLER_11_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_220 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_35_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_68_304 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_150_ VPWR VGND VPWR VGND uo_out[3] _257_/Q _151_/C _148_/B _148_/C _139_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_18_245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_279_ _279_/Q _284_/CLK _279_/D VPWR VGND VPWR VGND sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Right_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Right_52 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_55_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_202_ VPWR VGND VGND VPWR _202_/X _255_/Q _202_/B sky130_fd_sc_hd__or2_1
XFILLER_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_23_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_133_ VPWR VGND VGND VPWR _133_/A _161_/A _133_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_37_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_89 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_71_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_29_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_53_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_48_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_1_217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_49_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_360 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_49_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_252__20 VPWR VGND VPWR VGND _277_/CLK clkload1/A sky130_fd_sc_hd__inv_2
XFILLER_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_23_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_278_ VGND VPWR VGND VPWR uo_out[7] _278_/D _278_/CLK sky130_fd_sc_hd__dfxtp_4
XFILLER_5_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_52_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_70_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ VPWR VGND VGND VPWR _186_/Y hold18/X input4/X _203_/A1 _256_/D _200_/X sky130_fd_sc_hd__o221a_1
X_132_ VPWR VGND VGND VPWR _133_/B uo_out[6] _260_/Q sky130_fd_sc_hd__or2_1
XFILLER_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_78_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_709 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_69_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_0_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_236__4 VPWR VGND VPWR VGND _257_/CLK _285_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_75_233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_48_469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_63_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_66_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_92 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_9_329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_40_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_291 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_32_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
.ends

